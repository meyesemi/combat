module gw_gao(
    rx0_de,
    rx0_hsync,
    rx0_vsync,
    \rx0_b[7] ,
    \rx0_b[6] ,
    \rx0_b[5] ,
    \rx0_b[4] ,
    \rx0_b[3] ,
    \rx0_b[2] ,
    \rx0_b[1] ,
    \rx0_b[0] ,
    \rx0_g[7] ,
    \rx0_g[6] ,
    \rx0_g[5] ,
    \rx0_g[4] ,
    \rx0_g[3] ,
    \rx0_g[2] ,
    \rx0_g[1] ,
    \rx0_g[0] ,
    \rx0_r[7] ,
    \rx0_r[6] ,
    \rx0_r[5] ,
    \rx0_r[4] ,
    \rx0_r[3] ,
    \rx0_r[2] ,
    \rx0_r[1] ,
    \rx0_r[0] ,
    rx0_pclk,
    tms_pad_i,
    tck_pad_i,
    tdi_pad_i,
    tdo_pad_o
);

input rx0_de;
input rx0_hsync;
input rx0_vsync;
input \rx0_b[7] ;
input \rx0_b[6] ;
input \rx0_b[5] ;
input \rx0_b[4] ;
input \rx0_b[3] ;
input \rx0_b[2] ;
input \rx0_b[1] ;
input \rx0_b[0] ;
input \rx0_g[7] ;
input \rx0_g[6] ;
input \rx0_g[5] ;
input \rx0_g[4] ;
input \rx0_g[3] ;
input \rx0_g[2] ;
input \rx0_g[1] ;
input \rx0_g[0] ;
input \rx0_r[7] ;
input \rx0_r[6] ;
input \rx0_r[5] ;
input \rx0_r[4] ;
input \rx0_r[3] ;
input \rx0_r[2] ;
input \rx0_r[1] ;
input \rx0_r[0] ;
input rx0_pclk;
input tms_pad_i;
input tck_pad_i;
input tdi_pad_i;
output tdo_pad_o;

wire rx0_de;
wire rx0_hsync;
wire rx0_vsync;
wire \rx0_b[7] ;
wire \rx0_b[6] ;
wire \rx0_b[5] ;
wire \rx0_b[4] ;
wire \rx0_b[3] ;
wire \rx0_b[2] ;
wire \rx0_b[1] ;
wire \rx0_b[0] ;
wire \rx0_g[7] ;
wire \rx0_g[6] ;
wire \rx0_g[5] ;
wire \rx0_g[4] ;
wire \rx0_g[3] ;
wire \rx0_g[2] ;
wire \rx0_g[1] ;
wire \rx0_g[0] ;
wire \rx0_r[7] ;
wire \rx0_r[6] ;
wire \rx0_r[5] ;
wire \rx0_r[4] ;
wire \rx0_r[3] ;
wire \rx0_r[2] ;
wire \rx0_r[1] ;
wire \rx0_r[0] ;
wire rx0_pclk;
wire tms_pad_i;
wire tck_pad_i;
wire tdi_pad_i;
wire tdo_pad_o;
wire tms_i_c;
wire tck_i_c;
wire tdi_i_c;
wire tdo_o_c;
wire [9:0] control0;
wire gao_jtag_tck;
wire gao_jtag_reset;
wire run_test_idle_er1;
wire run_test_idle_er2;
wire shift_dr_capture_dr;
wire update_dr;
wire pause_dr;
wire enable_er1;
wire enable_er2;
wire gao_jtag_tdi;
wire tdo_er1;
wire tdo_er2;

IBUF tms_ibuf (
    .I(tms_pad_i),
    .O(tms_i_c)
);

IBUF tck_ibuf (
    .I(tck_pad_i),
    .O(tck_i_c)
);

IBUF tdi_ibuf (
    .I(tdi_pad_i),
    .O(tdi_i_c)
);

OBUF tdo_obuf (
    .I(tdo_o_c),
    .O(tdo_pad_o)
);

GW_JTAG  u_gw_jtag(
    .tms_pad_i(tms_i_c),
    .tck_pad_i(tck_i_c),
    .tdi_pad_i(tdi_i_c),
    .tdo_pad_o(tdo_o_c),
    .tck_o(gao_jtag_tck),
    .test_logic_reset_o(gao_jtag_reset),
    .run_test_idle_er1_o(run_test_idle_er1),
    .run_test_idle_er2_o(run_test_idle_er2),
    .shift_dr_capture_dr_o(shift_dr_capture_dr),
    .update_dr_o(update_dr),
    .pause_dr_o(pause_dr),
    .enable_er1_o(enable_er1),
    .enable_er2_o(enable_er2),
    .tdi_o(gao_jtag_tdi),
    .tdo_er1_i(tdo_er1),
    .tdo_er2_i(tdo_er2)
);

gw_con_top  u_icon_top(
    .tck_i(gao_jtag_tck),
    .tdi_i(gao_jtag_tdi),
    .tdo_o(tdo_er1),
    .rst_i(gao_jtag_reset),
    .control0(control0[9:0]),
    .enable_i(enable_er1),
    .shift_dr_capture_dr_i(shift_dr_capture_dr),
    .update_dr_i(update_dr)
);

ao_top_0  u_la0_top(
    .control(control0[9:0]),
    .trig0_i(rx0_de),
    .data_i({rx0_de,rx0_hsync,rx0_vsync,\rx0_b[7] ,\rx0_b[6] ,\rx0_b[5] ,\rx0_b[4] ,\rx0_b[3] ,\rx0_b[2] ,\rx0_b[1] ,\rx0_b[0] ,\rx0_g[7] ,\rx0_g[6] ,\rx0_g[5] ,\rx0_g[4] ,\rx0_g[3] ,\rx0_g[2] ,\rx0_g[1] ,\rx0_g[0] ,\rx0_r[7] ,\rx0_r[6] ,\rx0_r[5] ,\rx0_r[4] ,\rx0_r[3] ,\rx0_r[2] ,\rx0_r[1] ,\rx0_r[0] }),
    .clk_i(rx0_pclk)
);

endmodule
//
// Written by Synplify Pro 
// Product Version "P-2019.09G-Beta2"
// Program "Synplify Pro", Mapper "mapgw, Build 1530R"
// Fri Apr 10 15:59:35 2020
//
// Source file index table:
// Object locations will have the form <file>:<line>
// file 0 "\d:\gowin\gowin_v1.9.3.02beta\synplifypro\lib\generic\gw2a.v "
// file 1 "\d:\gowin\gowin_v1.9.3.02beta\synplifypro\lib\vlog\hypermods.v "
// file 2 "\d:\gowin\gowin_v1.9.3.02beta\synplifypro\lib\vlog\umr_capim.v "
// file 3 "\d:\gowin\gowin_v1.9.3.02beta\synplifypro\lib\vlog\scemi_objects.v "
// file 4 "\d:\gowin\gowin_v1.9.3.02beta\synplifypro\lib\vlog\scemi_pipes.svh "
// file 5 "\d:\proj\dk-video-gw2a18_dvirxtx\project\temp\gao\ao_control\gw_con_parameter.v "
// file 6 "\d:\proj\dk-video-gw2a18_dvirxtx\project\temp\gao\ao_control\gw_con_top_define.v "
// file 7 "\d:\gowin\gowin_v1.9.3.02beta\ide\data\ipcores\gao\gw_con\gw_con_top.v "
// file 8 "\d:\gowin\gowin_v1.9.3.02beta\synplifypro\lib\nlconst.dat "

`timescale 100 ps/100 ps
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="default"
`pragma protect author_info="default"
`pragma protect encrypt_agent="Synplify encryptP1735.pl"
`pragma protect encrypt_agent_info="Synplify encryptP1735.pl Version 1.1"

`pragma protect encoding=(enctype="base64", line_length=76, bytes=256)
`pragma protect key_keyowner="Synplicity"
`pragma protect key_keyname="SYNP05_001"
`pragma protect key_method="rsa"
`pragma protect key_block
nGQjNTRggZWOT6sWc6oyraDUFLfWAO/HbLF6wXbCqXPNp9WCDJpv1rHVczOIVgncR/b0+UeSwebZ
OxlPzCeuO1qPl8FPTKiUyycPd+J0aSTr5vl+//g43DlAnrAZWpp+9NwkyX7Tl4KQV38q+/ZFnqAd
fKrxDpwkhDu4v9GmdKTtVryneeZJtk+qfqQLeux8ui4DI7WokBCiLCcnunBZc7zPDJ4RNHhhj/d6
kphLiA+2e7BZhQi3+S17OFvZZeAZqB9QHyWn8tsgCw/p96pTPtatJ/h1TGMYgxgbBmCeWweLMmye
bCwg5pbhghYptD2zVIQFJWuiylXMfypQ3ZpFdA==

`pragma protect encoding=(enctype="base64", line_length=76, bytes=256)
`pragma protect key_keyowner="GoWin"
`pragma protect key_keyname="GoWin2016"
`pragma protect key_method="rsa"
`pragma protect key_block
x5gHfLwQ9h6IkqXYFQsKYOoMTbgAOviKZwc0Vf339pYT772gCzJCT3UDF+YsUsYbK+Pq7BKRT6Uf
HBulNYuf7y+Ku9k8h5gb4vT0dUa4DG8OSdHb7R0AC/h0AeBTlns2hBJ4OSQGxyyNBp2s9HonSdOM
8ZWZFAphVVtPxikUpfU8q9qzyHTb9jMLF3VfqHt1hy3qcsmu5t+UPmv9c2zjTl4NXRMUl5483dXo
fMq4baFS/ju/wiHFuRhteazMg0mM6BfGhtM2aDlFaVzlnFbwItgar6Mu4Fk1u80ynR+wqXfj4ur2
96zU62Pm3UBbG8dYUGOAgfAhYDkhAs6USGbytQ==

`pragma protect data_keyowner="default-ip-vendor"
`pragma protect data_keyname="default-ip-key"
`pragma protect data_method="aes128-cbc"
`pragma protect encoding=(enctype="base64", line_length=76, bytes=7104)
`pragma protect data_block
S64wz9lq30aLaC+kL/X10osfDUSymmrQf6hdQCYuLnmlW6w0Fzin4aO0g/WUobnGsoCOY7+vwaK7
shINCGen4o92p7HrSWBdN+5Baowett5dwKHQqJmKXDf8kRu2EUM6L5usvI7gmjwb0Oqr0AOxGdMA
IEt240OIHMHC5+4DWcK1R5uW4oisAZTZ0NJomTQDaMYTf0vbCXRvBfHpZ4l5DtYYykQ+1wrCdaX8
sSH+7Kja8QmLHvKxnpa8f5JIgVG/ucAiaLjJCwWMxb9Jgg651lo4it+/5Tpuo5y2qsnz4H1JMNUn
Uj2Wb4mlOEYAAuxfOQgISpA8CPBcEc7sbHGRaiqACMoKpmzuzNxNUD8P5cv6ovUqQfJUioqy8RZU
ncsdMPHyh5mNATv+rgnC5o/KV93EFFByE293XvqXEYEjt9+B0tjML3MngPfTex/cJ2bRYI1Y29hm
XTL62PjJKbMzmK9NpFeIkHzsZDbc2u2z/BIavl6tVtDLm+SAcnppavWyK/5wQreqZ2yB53u9z2o8
LprLjQ9sr4VB4syjJwQmDoIF3R2IbM/QcfbvefBq4dq5wIAzfUOIsG7ArZLpKq5bpD2Zb8A9OHiX
uvKXXGCAt2zRRcVLod4NupUa6X2EHnU26zdjJmoMtd40HPn4cS1oNYsj8oDgnMRuf/Usf2EPCPzZ
zBwI1jWvbx/LDqAKeiJy5p6Z3ppYHfexLl4KVFJwvZN/UAIWIEdE4gMnasijR0V/X7zNIff2Z+mg
Vst3itLdrWLhIpU72gmh+FTfXmgP5G0QzeUXu+8N1eSeRol7/A0ii/TmT6olTEgp5qz99PEILD9D
dwbTqx6rbR/vbvZYn5A6MKVaJHf1Cf2AGsVHwSde1kyO3hEKtQ4r9nRWUIdDLZuN0jDbKAOGjSOj
cKQrNjYtn3fCdAE+vAydqBHJo0aNdCmOVR4Q2pRU6nYrm/btQlG2q7hLFtC/KPp2DUkDmxN8r+5B
jtXBUi4kv0tFiBkb0PSxuTRWBbmxgMHvu2TByRH6BUq6yGS45JSdbjpP0iYwguTga9uQlQJseJvN
j15bPLNnu23qzXFj4YABLhVMn3u2NXCFJtuYMqFQMW1J4orX1gR/oDz9x64hSD6+sdyOMqp9gEDe
0WZRRJAd6GzrepdeVLDl8wkUL5q2LruU+iqjEWV6S9w6E/+nxR01/BtxYLYurB06WOIux2dQ288m
+GGE3sZDqGx+4Z8RhX1zXr+jWRREuhScq0o8HakXzrQJ5d6LY3XsmvevNbnVF62XHGOq0jtREcXU
H1rGoR5lC3ijAvpx7b8Nk6N9VmI+ia0y17PcS32wivatHlatOvDz21513YSpkq/Yw2A6uJRl8KVH
Jj+kLgnAtJuMsFxxnHHDEd0DwbhpHYNlklIcez4hcNHHcW8UY+129G8pPPfxT0aJwrvc8xdF3FO5
zGC7rZuAhq3x1cJ/zlTFsepDtjwvqoqUCODzgXBkdDzWftJn68ittbbm+zbQzXZHy39+5j/0bQGq
xrYRoc7uHFk9KdSbpbDJdvad2clSy0ty9w4csPYjbsz+kkb94vouUIdy2WpnMkdbST/cPwsGLpfj
udJD5z0gsk2qDLqeePnl3U/C9moYz+Cw5pa2tiYU0V8BmX7+oShtCNHaGx/694KY617H2GQzy3oA
m7axRdZFb0Wf5dz0Nx2TmDvYGlw8284EwrgIzrOmqP0aBAPXESpUujnN+olGWShGRd5EtgOyQLgI
HhCppZtOjMPSKULg1NinMUMFPFZIn3dNlRGv2wFaiFFWDgFJnKxRNHujBhtdwAf3yifrXHjvjlq+
rdBW/36IfXTsD2Hk9yW8sCyFEJ8thBI9kX8v9IynnWfRY77pExP+MXu6n1mMsAGI5+NMIIvtD3/I
8xOHQ4Fm3nw61qa/ENEbZE2xLwnNBdbKhRkOJ5E61hofSr+tdUO7JXbd6HEDKhyQgNHJRVAlCaZg
nxVNBSyNe05LUxwkXsArTwvBn8XteTvnwreP7Rvd46oUPX9at5gkj45CfbJkoid5ejxoP7oRA8pc
b+LtAJCrMLquvMjrcRKEjqw+yyUwIcTu2KqmtaORXZbFfDMTQidCAL5iiZiQBMmtRO3/2JWSeO/z
yisWQmRAJxgLaoyfQTxLqqv183VR0dQI10GRQNDUNkuSEADQyOOj93ejJfRl7bMQft7oV6nVSCuQ
y4cjRGk4zWKW0i3x9RhGpv3MBr3PSrgrf0dmtM+SQAyshs8XMHzJevWf/0Y+78vbIDJJg1KwCgc5
uDOLVwDKf4yKpJU7loF9aKfWzRojoC/RpzyT9A68n5qc+QDWvPhUBWhrKN8weI5h0z8dGcwY+9z9
yED1Ockg4xGHaqcWGGWbPa5C1rZUCPgFkHsmyLX8W66yGl24nohnk0O/GNwCNhNzhVwQwtkawho2
o4AiWfYhdFKXouZ/racJoqYuoAV/t9cIMNZEG2q8vvHIXNf6/NB3QDyyNrxBmJYSwEABPH7rCvDI
rDzMLY7dGRZ1CgyuP2Ge2RY28vqO1sN05e4EbXxxz2GQTnvAf62+oTQg4B3cMKNkFUzO4xLyV4M4
A3r8mmGj/Kw5MHLbs8dl44f+P9vU/+N7IiQWRgPdfhrNIPYmrRRw0o3UEl5GQMa7ersm2H20+i3Y
FLw9medsYw903pVmzIBH2R1YUdNrYOquqVdI3cEjOHbVLruEmC9CEP6s8mRyi9ixwNK1ZGF7StYb
lYUvkpMh/FbEOutMh2dAYwuCQaKcUtQmP3d/SMDOgrDKXiJKqE6tzq7W5TDy5HWT/Y43/TdUF8BK
0jJX/krAu+lIqq+KfAkrBVy1aZR7TVrpuJptvSWUogS/ZKOQecBI+DScbiM3p7ZHod5X9Hlt+on0
Eix/WyX6Xh7Qr5AqZcNwvF6rTmcIBKjZv6j+y2Flnb7VMqDsTB8bAOoBRPnWW7yEWyy4GXrxoX8F
Pj4hlK/sGSmfTI1ioE/HOfBGFUrMTCaxpq3uOcMxBQeeNoZJzL1HfxDFntp0z1s/Rv/KJcGluUaU
LRAaH/I5r9XgOinwSRcjpBrxjS+uiwZXJu1JuCQz+pQcsbsP1hc1ZM12XHKr/G9/xkPgzCiMVkLk
E0wlaFyCxuwgxb889oZCDYq+huWYcNbgMGyi0aW+QYuE8Ha9YlNJf3A3XJxk8tTaxhWqXNp4THVn
ZU7UM9mZwAvK6ef4+/UugG5R0gLQMPPSa4+TeXQDgSYeCOWKs8fwhKrEpzgFgoPv1e20fd7MS/bU
Op1AIbsXYQcxcPvkx9+QPszLjD2V5z1vmt91ndI0sgzflNwbUVdkhMwrBYowMnJKdCru7q6mqi/a
mCV3l5rBjDVHh0LiICc4jMrrSo6EiLhNwWFJWowZWTCkUNIZNUKegYjpBs7gmpuwndeGNxVfXCZn
iVlTRNTIfWj2fb8GIQ/mJDa7hzFxv/21KhESvnTDuaEjy9HaxR0+OljsYi6owDKtW/cj4ei5Khnn
kKXigqdMoPQnBBy5+Dlu8xs2AWSIQa1wUyoGqjBATErO6LXslghIbgq3y3ExZTY5kf7IKKLBmQaz
YxJh3X/LJLQkgk7ePJveOrVRNEA1BMm4TdqAFj4pBlAUeMcilNPhQ+gX38QGT480Pc2RFSWW1+ZN
oefjAnTTwBcZ8z5Yac/0qMttIH0mDph96GRuSx8VEpQ0hr5VAkTVoUohABBRUHcb9Ls90mRafwUA
lbI3mwbhRsCkcsDJB4jutp3wOCt0BVnc3b2+PBN7AjQRSASl93ofLhAxfVQ03l1nSibvSWe1+wbG
2dUJy5u2M55OD1N5tEIcI6o95cLbNOx36bQSpDSigg8keHtqgKYe+fFnQZUWWXohOI5mATn5hRPV
KiZfXbB31Oa5A3DDm+jb5C4+D6mSI2LLcQZe6yknElDChlD9GQhlBTqUAG8cGVwlMftOZ5E8BwPe
rkBZP4Ih+w5WxPnkeYmydhqWLnoSSI6HIFK+gkJzsuTlBOU93wYBBG6Umg67l3bAjI4Xib3N5jiB
ZbFxokxItCnNtf1FFaLK0+2KHPTAPbuhOE2o2IYQpnab8Zegs05TYPyRSf2/7WpTtkDdiF7ejKlc
sPA+xM8N6R6Yrwakae3dS+Mu2Y6OntbT4U51BJmslkUEf0mWTY96RF1BVKUL5SVRgCqHRAeMyHaz
qHvSApD1czKbgf4i6g3q68umeUXAJJLiegmNd+yLjbdIGrlofjvBhlw3n6umwbU2Sqxw0NQM8HQ5
K6XxvdnDQ1OBfko4XHIFhhkhse8agYli7HJ0cpOsC0vaeHoA+BTC0lAKOkOLLD9Q+wI5y2lOBRUI
R/+2kC8ndhlEWoROS1M+bMQ8AURisonhvfmHAt62wu6CSGlbYwkp1I3sUxtx9kMmPnGSe5NHe1Jr
wGSchJ1g/D0weviUf/8UAtojoJiQUi/eezHzww2DQfz5PvREUkVQC1Se72W8wF2L4ATqFFaua12b
wGFTzC1JLsaMMaPmL8v5S0d4vhhorHtY4uzrMjEeS8uzcjyssxaVOE/ZLklT7bX8DKdlmIhWRAKV
qHHvdKv7weZ9yTsxXKWZaUpg4MHP0v0gdGecJ8xkSageBrXGZp1pI47y6W0v7bc3EMyt7rV7D2nM
hwUGuqQhktdwoQiLapiHCtuLi1cKGeScbabmqW0gFXV5ooMTafetu2mHFAhx6q02YZAPQhfcosP/
gwCqIcK1YPBEyJ60SkW9/KGp/K4XCOuyqgbcI4RHUPXCHgI8cVy2pRTbCRMb2mi3xA/Z90FEU3Xj
uQrcGrPom8pyR5E+2+9LpynAldtSRq8Zcv5RDP9JX5UzC46Wz96g6N+mgtkn2HEf65hkGMeE4lHl
7QkSgTEPQU95gFeFdkSbRIzkbBuFoYeLSRg+C2NVZafssUKr+hmVdhlxpaBI8H/Pm8bhBdMuTDXe
baF4PjmAlt+jvXOW//65RpWxZIA7UMjfPM0qvzyqNa1pxutYSAlv2o1PcmRbP4FWJgREZrqHDODh
tH6WmdjzAX/aekH+OByWGjNbusM18D6S4LlsGX3TIzolLYTrISa2x6rD/dhMH42XZ3f4Euhx3p81
JBGaLYR0T6RDiPaxX6lS3M5S/iCG33e7TN4pN6sgdSsnC1dGZG+R0hxlKTJ8/uV4NNtzkPA/n3Zb
V/Ygx3XbsyC5jh+IHQvpMLdvbbZi3eiwvHwY5FHbhbBG5/UA8B1WTNIozV+Inb6mH6Ql6upBbU7n
1BfBMCH3b7kgLpqj8FycR6TbdsifLKegykv4rvvIUfrFos4NRkDaZigtCaiIZnVXVpTO1pWb4zif
EgNlCkNstuHrqcoEPD3crhgsmeH6Xf/rz8L/q1j9Kgqpq9qPUwUmttjr3ADtq4sTp8OgyDp2JaY4
6vYD3iIlvsrZsntzpWMm6c9TPsd5cTVpBnUWd7aB7v0eMN8BEbrJcwZPQef53ogY0XqPYaEL+gko
csex+bKwfWUBCIa0CQFsVSMTJe9XfCiItiSDI5COuXus8rISVFLgwl9d8kiYz0wW4Uc5/jGhwGVX
zhQTdRp0cN9HA57fWmind5vjXwI0qe9yRK78v1upOq1Vmms4KMz/teObjCkPbX2B9HaUQiRhVt33
tNliZfjsVNVTY/oHA5nCz++NA1vN4U0qKQhI2MagqKVuWvCmdyqLP+lf8FTnYwrGXYeg4MOZ0T0T
WzhUhv2C/dNmk8N6/bBUkJuH+WXhb1pveUkLBM3M3YQIYKbjMZTNooiG8dvzTIWbZRipW0rfltGg
rxX98Xl4nw43GXLStEFK8zFBjSoYFqVRMrxgyT+1VKGR8kEYIam3L1ZeP2qWvw7+Yv6+8rFZzKeZ
fVjENVwZ+10eIBH9pHtOZtC8NMv9St1efR33q84L3UZ9YoN+brKClkspTGiw7xM6WMZxur4Xj5K7
3Ct95Si7wTDo7hrfsHA7EZhyCAu3CDJg30Yc8iHhD6oCXL5Jbn4cgi0JAiiIUmXu0lXra4o1OrJG
OEmhCcpHIaRtlsDuyhat8zQI33wGe7LmOThpLb65qT3WWK5DJVxnJb+BNALWwz0bNckMVcWjPjvZ
wbWRKCo3RJNQXFiYWGpDlujc/LoTckBnG42+9RtV5FteQdb3k2KWxs+EyDzmWuwJzt9tmff0eZZC
gktiPz3lhmWywZtI/GZY4E7D6zOo8f/Gou79Sll1LmKjrJoYerB7+BHDEkWr6bl+uR6LvuCO1NMh
8G/+IcsgDLbpZB5T0XfebVnp9EkfVSklT21oxBixgi3KSFOi9eWAJp3zXrTY4RlxpBXcMTr3gvlF
chOj9VsyNQAX9jp8eIZrx8UAZf0uBe5I9WVQ0cOGJDdwumtgdvmAwYyiHwzyGNZ0lUMkzKNMQtXA
2Gf0xVP0mkRcezCmiqoFTGu35veszVCnM+LYQe9Vf18LaD4Cv2ztI1+RjTTn996RNBHkUR0n1ZVR
/JOkPTQGZ2I7wRc+UDlZlZgbyPSSfBJJjoDBUuNGacDYSB5RMhrmKwpu4ej7ESSqnx9xiLQRCJ8k
mhlxgHN0L4RyNYLHfuQNU12gepUGGjy8CgrLxeV3SRDIRuWqMADgfDgLrypwBqPorM2sMs9ptX68
ktZFXcwxJdcqo7diINqZGmGrlEIfuh4cTGp2j0BMfMgzbeYUpfaMOC90U66LKoub+dp7aaBdyyzX
OSl858zl6Lw6wD+bMtiqGboc18KwIF7NyesiOte1SF1CjCbIawvMNlAO7ORmQ5RZyOUKgnkOiTBO
3vgakwZXogeXnYrZXjwAKHlPuWAmiiXRs1sBu+slXY6MDMQv5sp6AAd4wj5DD47Ekvqa49Im77Pl
NnCFOod0mtE0+999pgisGX3rlFq1CqsapTgnX4XvsCrYQmxZsdAdIbjiQxIWZZGwy6zAFPi/YY5+
l9MTHXZBO8G1+iJtEENsF/RXb2fdkDj/p/VhmljDFL5DsGk7Iuk+X8OrazniOoDPqXtFaPPSb8d7
o5CwXbtQMmuthC+kjoomZmrJ7SmFneiw9p39ckPoZA2RqgYsWYTMD0wcwAsTHe8T32VGjAxHXb4w
vTIAVNH5wpxDKNOAodjFMSwz3qBcghDJwctosIPna1U3oU6paurBSDH1fPESGHShTsuCDPkNt/3A
ymgFnsOCYBzu6zuo/jECemOIMVLykEINTED/91fxnmmgmX0J0flYvVtq4MNZ7qWX/Wo5ssrMIMkz
+US0P2+t56X9yc9EsClGzRzNJdSAzFM6c2jZIz+p/VjrgKuyT0lhQPWEw9G2WUpB4xTtPhTsjQ6v
mG8o48RabcM9zOjLqYSQR87B9BHH2pD9pf5QtXTDjkGO/b6++aycn4oNCN+v+vrgGJAEHC2N13cW
RRh+i/1eIU5DUwBhFf5WegUCuhV5e1aNoLzmgAGOTf1evg5y7IJfTgg0FsnHXgMwBEYgCtiAEjLe
0+Fs1Yd0yMMl4q3DKH7wVIpZQBeYYVM+ENr8w9U8jS8N6q0JPGSbCNA3GQaqtZvsL4+RiJrXe3xr
vUIoMnxkHHR+ix3y/23R8hvVvhnvOnx/0YIB0fBy/ema0AnH+iBSjFaYLM7vuJvyCr4Q769jzT5q
u7RGBNQo8mXXoFmEe/suMcTSbeSuK/hwYB12bAyIDoaLToVOhHryyR514+pQCMz5KgS66TV9D3oi
a/3e6C0Og1t4KWg6it+TGLGw8RGJPh0MXoqR7y01no2Rpjs7MzlLH3E3IYZambc9YpdbtDCasv8W
Q5wKK2d9xr7MAU9XOTwscE4Xv9d6cr/bfirH7Lvjg2LWz6KWEu/UAn0YQZ+V/J4VsTn/bVrk/eaX
PZpSsFSesf7JBcYVGbKbmSTCH9iYA3dW//LvyPXuTz5V3686tABQqe521AR3OcVGr/2VHkbt1upz
PvROv6o6kNCj7NZTUGGkn4ZIjnqqhPuDPqHlVtHGN3t0V02WlcB9gqiVB7Z2sGteiBHKp/yEXja4
WbAWTDyJ7DqA36BuJwDo3vAQFDA8/dAvepjqYD5r5VqbJqudRyjsHuOLEKbdtJGZm5zWvGYYoNw0
ARqR4aiIMMSp6nIJUdiKc0lWZuie+ubOIBGZoX6OjWbm6NGTODFAD61hWGFgoR9yL7yhLuMtcrGg
1TKst12FTuVTDpT519TrwCAavJu5jLB6vVooDxUWfZRhgJOub7NYxx2A4aj95j5s8TuFqqdLPP0T
H41qe26XL2EUnRsQDXFX/JkHH/mNpXkNxNqJz/c7h08UTGn0tsEMypIkGYBirhZWkRC6YBrKAjzJ
NkVXRmNFKCPFwh7DsIYwq0hUjS6fd5KB4Sh0Go2a7t9nBhMVMr5R9QHyQr/CGMKLzvgpaxXTpHR0
mTkHjJNAeWzNVdYzTWG3sLqhC/9dFOfU6F3FLuN3WlsEkpyv1vPQ9iGl3MND2k5O3dPIxobPRmf3
o0T1oRw3gEQ1Kj8777jZO9I8Uny3h5KOv7pbKlOWeCjWb6MJ6N4Ct0TDBq++Skyv6YJipDIhJKqa
pL9IgvVUPM9ZtveUpCFTSnLh9WPRuJOTkQoYQkSpyPQuk0z06SOUgBU0Oasif2RC0ZOhOUlalUQ8
iWlh08Dv79eNGZIHJ2wstW67cX6d2mOR1u8UerxZXwuOWv9t/tKoUYlGruZ3JQ1LwWVlk4y2K7/E
cXY9I9YCQPJrMV7+Us2RifXM900SRft/vmFecRAQ2L1Fw9cy3hd7YRBcUpf7fL5s3i0a11xQQxXB
fKiiV+Dg9Xj3a7HX/u0bcnQ2VDgemdvOJMw2cNl/Q5S6zTYjGpvaHwFCd/46YWACiRCG/5cKoN/N
ueBzxbkXfVAkf9VJNTy85ep1a+NzjfuaU58ahtvTO9miRK2ZbucCsOeak61+6CIbB2es45bLzRml
6xUZSEsRZDN3t+uvmw/ujPADTmMzltXFpRqu1MmSaudaOK2aDXAZJj4/t1SdaNwAi4rMr64MWCvM
8GSpZVXHAaQ9MRoomQALFHzCNXBftQALac4Vm154Rr9JdfpO+C2zRAS2zrv0jBukrxc+kjOwKyJ7
oAKfYroPTvkgcIknimdNFqohPzHvcSroA3qsC5aJ7jnQEYtqbko+0p+U6cC1i/x7G72SPOr2cWep
jMkU1vNJv7a30OSBx4zak5x6FN78jTeGb4CUaxVMBVHzpYdqllvYP+7PDZeZ8IJcJb9VHzWWL+Vy
SvQBtEM4uwrUSG6Bo8Ecj3HBEktuN33NYSeSPXzzuMySZdAALD6Es2xXigIVqPCQceUDCVOe3BlK
WHF5B9WHHOL1SmhGO2VBaGYunZCbeQdtI5p0jnTVH8yXQHq4WzNk/v+igL4NWTOOs4Mp/prj+wkE
BCttwh96l3EqP2y27GcHnn6z4FYKMueLuhDDh4vSVAReMFkyObjkr958tFwKukAg05mM3Pgh/LmX
3PzsF4PQXOQizNvIyNLkHZ3B6iWi8rtPs4KQKEu5ZOsbQC+9
`pragma protect end_protected
//
// Written by Synplify Pro 
// Product Version "P-2019.09G-Beta2"
// Program "Synplify Pro", Mapper "mapgw, Build 1530R"
// Fri Apr 10 15:59:50 2020
//
// Source file index table:
// Object locations will have the form <file>:<line>
// file 0 "\d:\gowin\gowin_v1.9.3.02beta\synplifypro\lib\generic\gw2a.v "
// file 1 "\d:\gowin\gowin_v1.9.3.02beta\synplifypro\lib\vlog\hypermods.v "
// file 2 "\d:\gowin\gowin_v1.9.3.02beta\synplifypro\lib\vlog\umr_capim.v "
// file 3 "\d:\gowin\gowin_v1.9.3.02beta\synplifypro\lib\vlog\scemi_objects.v "
// file 4 "\d:\gowin\gowin_v1.9.3.02beta\synplifypro\lib\vlog\scemi_pipes.svh "
// file 5 "\d:\proj\dk-video-gw2a18_dvirxtx\project\temp\gao\ao_0\gw_ao_parameter.v "
// file 6 "\d:\proj\dk-video-gw2a18_dvirxtx\project\temp\gao\ao_0\gw_ao_top_define.v "
// file 7 "\d:\proj\dk-video-gw2a18_dvirxtx\project\temp\gao\ao_0\gw_ao_expression.v "
// file 8 "\d:\gowin\gowin_v1.9.3.02beta\ide\data\ipcores\gao\gw_ao_0\gw_ao_crc32.v "
// file 9 "\d:\gowin\gowin_v1.9.3.02beta\ide\data\ipcores\gao\gw_ao_0\gw_ao_define.v "
// file 10 "\d:\gowin\gowin_v1.9.3.02beta\ide\data\ipcores\gao\gw_ao_0\gw_ao_match.v "
// file 11 "\d:\gowin\gowin_v1.9.3.02beta\ide\data\ipcores\gao\gw_ao_0\gw_ao_mem_ctrl.v "
// file 12 "\d:\gowin\gowin_v1.9.3.02beta\ide\data\ipcores\gao\gw_ao_0\gw_ao_top.v "
// file 13 "\d:\gowin\gowin_v1.9.3.02beta\synplifypro\lib\nlconst.dat "

`timescale 100 ps/100 ps
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="default"
`pragma protect author_info="default"
`pragma protect encrypt_agent="Synplify encryptP1735.pl"
`pragma protect encrypt_agent_info="Synplify encryptP1735.pl Version 1.1"

`pragma protect encoding=(enctype="base64", line_length=76, bytes=256)
`pragma protect key_keyowner="Synplicity"
`pragma protect key_keyname="SYNP05_001"
`pragma protect key_method="rsa"
`pragma protect key_block
DI4rXVSqQQakdxUiFbNMpUcFqLtxiH/v9VC2fotO6RT5oJx4ujfd+d8ntglwi9SznfUhuCDdANfH
XYMgV7tqilOQ2ZawjyjFzCrZ5SPXrGgsruT0nRljnPbi6qkiFtugOcQTRLawx9T7//cBM+KloXTA
NW5UEesUVY6XIevfIUZGJ1ure5Ny3juAG8DwrfgVKoVsVbpFHGqkn14/CuCrPfgd3cNIeMnz2tdU
fIIQcJuw7/y7oxsPIHnSNjduB2VlABUbTul3/U+MLlIz6QrQXnGGd0gsk0VzmjNw5t92AUKNXFJQ
KgZfLCLpjgQ/ZbGsMSNTxIFdLQdlxHMJmC0vaQ==

`pragma protect encoding=(enctype="base64", line_length=76, bytes=256)
`pragma protect key_keyowner="GoWin"
`pragma protect key_keyname="GoWin2016"
`pragma protect key_method="rsa"
`pragma protect key_block
BJq830S/kOcQBA2JJ2q4S6I8jB9jjQ+2w4M1vD4Tqw23sKPDOhifxjr0/o3W8kskkjrPH5ExmJnx
4+Ax8NsC3/y94RfnMYtaR48dVDd/uZPC+H97z8xQbMlRtAPIPBxmvbm2XF9esKwvNQk33qXslMT6
Af5S+VRtkbzP466p8XNJQwyztsU9oaM7FXV1jV3HosbJuRzcKVPEOmo4Dn/DOSxaP8rd5LPjoLqS
+itgiiOB0/sBM3oF4lMqNh90Lt7h7dN75Xc5z0AOiCtIi7ReGbnoPIxpLrTX3YY2f7/TaNJjwe2m
A2muDv33kmPJYj0Qn1mVE7WUxAUWY5au4KLJvA==

`pragma protect data_keyowner="default-ip-vendor"
`pragma protect data_keyname="default-ip-key"
`pragma protect data_method="aes128-cbc"
`pragma protect encoding=(enctype="base64", line_length=76, bytes=6624)
`pragma protect data_block
3l2m8UONmp/7H9fdVZbpxpmXcLOYUQ8E9OKnRpvBGbip6rCsDFnR2pm3cO97w6vSEQUEedB/p6Aj
/h2mgHyKH55lQd/cl26XFevQ9R2aFTRa0XsE16iM3l+26l9zxgiXW1bp3V8Cm1lwJrCXlb9g8csz
MicaRCchmotqO3GONnkx3CbxEXuTRUiCzvaJ+HR32pbbSyeIRE+9QoKHf+SvpUjiiLOKVDKfN+yO
V/hlP/JRcBFj+caIm2xyKPOE6BVzDV7GMN3Gzp/tXETSpn2VJPYO/kfffjJatoN9KUrNkDyCdiqO
mTC7HIHaF8r0LV1ARwFZTVLgsMfsA6LEn2Y72gNdrov5TkjzBEo6v7qP6wt7HB2lKdnadzorXLmd
HkTfdhXzp654VymWOfTKBBjqBOptswno278U17j3BsCY2MrDAYvEFiBFiLsY0QMhStKBao5Zh713
ydqixb1mfAJ+phTMuEGOQ65i0EznH6ZufSwRkFr8VGmK8C91VY7mpfcXa8+PCjxBb3q6QRBuRm+C
3Hx2j7U0tOUNrJRHVrHF4eAgRW7HNjWJKKHbUeIcy4WDWQn0pIL636rV5LKHFihL/JBR1Sfkl/An
UX+lvNQZC58NWXZzmwIixZ7M9J3YojVgax6pAcmLCEeeBb3fupFvdd6nuZ82cBkO+8bD5YS+S2dX
UgVxxne3j3fOaFLFG6xJgUn4tE4f05yzyhdmzbmR0RfPJUp6wGPVpjPBZUe+pJLBqkyMZy2BKeNi
NqiyBmwyVnsVyX5hijJF7ADFVMorhxykG7pPCtBzwyvG/vjGhzWDRgu6ygNJSduyOaxjGyHYe4kX
6zc62NCaCNCM+TYU6IFOHAHQAqykBPqxWo1sO7qdUQ6aSVZCJBlHbcMXEySMeyrd2v6JKDLob2Go
sCYaa/UgeOGV24GohLzOZf6Q+pfwsk1sOLh/fKG3pTRicaBexUlxKGK/nEOiD01Ui0E2FPxCPPAz
8m9MvNhS4YypRjqaaXPp/rCvVTdH6R2Yc8mib5sWGheA+bEC5/4uNQaNFl+TnIi8Uv67t11sitCL
dBIpSJAE20UKoqOIyFj7zBWb9EY8sg8sq5kKpX69S15VzqiVbmJW05lQ37PYTzBx9uClOFJtQz3p
PwK9ElVJjyXEGYBkCoA1W/s2XK4l9P2e7+r4vt0++ESgDhz1NG4PySpDH9ZyFaS1WNnAHai8QuqL
R0ZfVrAWTgnZs2v42bXpFTYNKAFtKJUX1+M8RXv6gxCqCIYZMTaSD14JWscky6a+vut/OhCjpEhN
buRMjvKWZyL3+i48ZbJ1hZbFCelA6NtYLqLLJlfQTrhiF/belbLcwobuzUYEOdhRn8tLC9nvYIAD
PT4QJnwbJNQSXUYGRSs88CbQoUb+9wlcy9VBvPHXY/Hb5t0ZJwPHD4uiv6UFQqa0ofkcei3i85pB
kh57JZpTV874fDpvtDuNawXptPNWWKfnnNm7O1Nn+SktFvNFhuPZ2YMSkGvuE8dFUn0jq2wVIGaz
jm3WZvJw1LaGAYXIbOw7SDfCsUGWPcxw7Lh/oGuxyjjDB+VtJKedwroHlcw9anSO/yHbVSCrIdbA
AiAzonjIrVH2hOW4g0KxkApos1pqUX9IDAdpWbUggcE110cGx4ICua+67OpSa500u+TCsld4W9sK
WqMv87AZ2+YTgyhUqEPrc5UcjXedR2sNw09QXnpGG1LIlSVtJmQFeNLaPVk7iFtbazs43Knq8M6u
AurQTo9ZqSzTv/be78JAt9jb0P89+tNWJo7YGGSH1DNoZgBTLXBbR0bS/jy2KdaQk4bvf8tp70oF
3mguU0aSEgcKmDnMteKjlLLZ3gAR4OCGj2jFL3TVPL6XoYcv0jZE5zlcDK1d68IDRKZQ9+LV/uwQ
CMTfouoibOV8oAWWDjCkgJ+TFfyFpNq0YEp2tRFTo75425VpJWNo9bBNoLXqcqTMZnLct/sQenEM
R6XvDPBVJwLKz59J/kCE4GU6EAJ6qe0FWMTF9zevxVR2l1R46AGvgfN/voYqQeCsYOr8Rkrnj+zk
4iKKhb59iHmFKS+uZ+help94/aug15VkD1Ooc7uQlgkn0ycKoCYJJFYvPatJZme34J9GMX/wMd5X
kWlCDcvg86brGMErDplRFu5y/KauEr5+nu5eP7IYErIAdyO4cFarWtz2F4/LkmBiQneBsbdUrv2J
mgbsTxb89hlcTRbJ94dgnFMbecDGabarmYqBaW8z7fO2nIWDpifA8D3lZZ5lomUiTwWF1mhWWPYs
aahMkOncrumq47svX6lljlIaw6OY9mIHOi9wVU373Ndv7wZelFGmlGw1Bk1iVeko5WEaa0Jh18PW
FLKfYzvpGBXz2/5Qpcvzexpc3X1l+/2m5O0Ay7LHiRDRERNFUehFPJDsNJQ3M515Cgr0OlpfZ2z4
NULHMFCwcajCxVZoA1msZEE42E32UaRsemG44o57vWq1oQAlRa2uOr45lkmRom2koFzOSA1P2m7L
OCadmVel85S3FVBkUqVSV/k330B7DUPGzDsRRvP9IpPfP5N9w2CnfGCqrCOKbaHzu1fePrv9wyCk
QNVY2HBcYwhtQRhUQ/dU7cR3B5/PFDvyRuV2jKDDgF+89lY+1eTbCJcGomelrpuC/1OuDM5Tk/A6
VLpOKwZhfS7da8j3baPopsZFfx1gQ54etbtJX0PhFBJWc/I9vmhrEzwai79QlxH+DAScXlvgt1Fn
MUBxovMgFFPalUwHpPZEVXE4O5b5In7smBEa1PEUiio+oqpNVyyA/AlTgkrh61KhorjrZD2tzFsk
pJCwhuomk+DyeYfQ7f/aMmjqfDhzJxgdD184kXlz50i7U7oI5sQaWpganaaOZ/uBNJenMugElHT5
Tpj3hUMC6KQY4PK+ZtFD34jRzFwXRjCKbK2LY2fhngtk0kyMlQ2/7tQUct5DD7CkJwEHbS/B982g
qcFrcKp8+Tyaw//zZTWZvzSw2WRDf+m5j6stEPieUz59tLOS98hEIwn6i1mA1lRU5DE6vGBXLpjT
LiYXIymwWiEx0OJBRdGCZmApN6z4SotZ1yjHZ4Maxzes902Nv5FGVgbnRDr/uEQflwbXL37Nh6Cz
+cy59a4ZyDSSwK/4MtzcIzyTC1XVWrPK+fffGml1QK11LNKRUb/FwcdFft2kxsG+QLk02YH7FlHp
Vkl9VM7AlSLjfS5N10JK1myGDU4z6oS8zfzIKLDKgyQwFXpksxI3W063jBLolqC0I/af/29KJdoB
y9Ir1jKTJaj0V0DObrsX5sflpV99Ums7ybvxJVJZAy7j493IT5VqYxK/UQbor0wRl7OjzUqxV871
hrB/DWI7MUX6Fyv9zbtH0/e6Jwsu23yLVcQthOW5aDkEyte6HOzt9dm1H7WFyMI8Uyj43W7yyjKn
S59Hq+xsxwC36sN9y0Jvkl1GcN9czMn5Exz5rWUdOMADMwRhfbN5KQvi+DTc9Ie9b7fByDHd4XZm
9Up69lhTB5SrTkvkzXgTF83Uw5L4uHck9fNWjaxdNKPYYRC6/vV2Xf0b00ldkUzJ+6jSCH3WR2bN
ywS9miudWx+PyVWZQ3OEkTSUFL9DWwdQqiiNwyLYZDqTkdhjTK1MRH5JOt87a6hwNApDWkyDzd14
bHWhg0u0tvoxjl621e+SmNXySgQtLTHywxGTAYQwNZGZSVnVoJV+LFm7MGn3Uk70RVu8Mr8BPTSe
k8IIDzoBWa0QhyT1+ZpHtQcDRaH1470hhOnZ5C1VXR/BNpJcNyqSU9Bvg7/W7sM9VhfH1jDK3stQ
v4jUOi1KzB1jWFsmEbXvI3kLWvxeHML8Glqkepd1jwoKjDjsN/yGuuGdtIPJm0j6o0/F/cbTAH/u
G8wVi/eMCqlI4C/MgA6nR3yhNlMZDPPbq95ryxQxKm0I/CDHPXE6/Nt62OGgaxZzNO8aDl339ojt
Ah0zfTTZCkQzoD0s/v0p7XdI6Nq28VmL9zGsTHsX4bA+QL66ydN/LXK9kO2LvBPXFbXwFWjuQZJ0
8aq6taMYj1Am2kdYJlnQw7F1rJ6cl9NwyJDxxvkyhCp4o+oX6K883r5U8DVSogf8tDUdCceCq0nX
rn3NRu9JiBsuYO84/oCvKqnHmLJpgtSCyYJWg3nSWSemsig2yiWTYsS4LvfrxR5oggAaVWoIHMu4
1+ZyFE/+sSc1uTp43HS0/2FH5dyhNCJ9WEwpk1JZdkoyk5Lu8z6TR9zKyJfdejCpKGuuO7aozUuk
Sxa8/DHyIPWd+SedZKNwiu6qPg7svBoZIoSq2c/Q1NrrYXGvaZm7YQXntwrjjf/0dbVYEeTj6KPu
BLKJ+gfidQZbhBfHUzGEwM3SBP0/qM69+JDYF2DSVlL+ygQLL6rQTACL4cwmjzNVG+ioA6J2FJJ6
UPPqtXblOXoHGspq3iCikm2RSbb8Vdi+9peP6bB8k2h3KLAP2IYdztlGglsP8bq7fcL4bmWkPFKR
aDB0FGH3bQPiK60aJ3fVbY6/Rm0Vsl1hrnNmhjYxX0J9cjz1R+J0dbp4VlmkdA2TFFxQARTfn+fK
NXCQKIIw4CGifPKiG1mPZ+YgK2Tw5ZlZopz2B47Gs2UMK1fS4RT3CxmOcM2ygT0uMUvRuDAx7x/S
P/6eVs9lcl9gMP9CRt++h6SvV9EF50F79RMtqEcUX8tL88CfknU7RTR20e/aVkmXTDUY9UND63Z4
29kQVtT7fi9yZT3RSDkzfc7s2aefM4VGEmWAapvpMGD22fULxYRBRmPUDrqjTknFBXmOD0voBBD8
8EYN5+p1qDkm0jqVEzX1nE71TEQymbQwgDPcd+kmlI/2qT4wHX4RB8XAX4SccwfTTDjqFdsNmpfR
sYKA/bsxlGiadZ3iNjTuPSX+s0rt1Av0SBuFQ+kwPt8k1mBDcqRys+GYYemjiCGkLLblHQDtoAfx
MAYWoI1oxYR4xgZMhNz/k9Got6edY0IKtPnw1N0FmMarkint0odXbyKrm/JvEEd5oUdljtsxZOS4
f5U2mDnnKtnT7bd83G4zjrHnw+or1h89cGmO9dwt2BfAphrjIwmF0nu3q5dQl9fVKu2fxPRLZnzQ
5RdRoI5mEk8w3FXpAbfqc92ZsZ2+XkEjqbrd9Bd9vztItaagxUudgoxIeLL5dbRJcnp5KxTB4757
s0UgQZrwzX4kbL5m7109RtlGoYZHpLjyJfp59FyDp/kBTf3ZnHWViw0UL8GlU6RhfpTy1FrptIse
jLhyF3a5ytlraoswxywcVm7TgDZQ4wxhzFebXOmoHHotVUwGd/IxnxRm0hHvcl36QAkDWCUVFFJc
Yo56GchDMI09JyhTodrrAKjm2r5PnRNzBSNWNdZqzTKfqsOzEvvVDOMU0tUGelgEl8C/7u5ifxpM
GZ/dfec4yVKhCDPFGqdrCD4TkYxmdy6GaxPyCzIbnLPEDDytM3YieVRPSCu8E3Z4AgijdpvNQvRD
zXPRarFRWPrxzfSH160hzVfOgk9HCtJXN8e7I5AdoqNg+dYiVBKfbQdSGOGgcXLxjOMW6t0fpiNM
I60DyYIKnE8Zxhxuw1juZGJQWGZG9Eg5mT09d6VFX5YGqr8x865b327UDLn465HhtNB6r/umAUTh
yjwsizp2wH7H/2hWK9saXCSZ/c3g2oWn9ty34NhtU3alKvv/GApCtpu9O5vOmyU7t8DCLZyZyyx2
vPdDHJ5YScJeQmcN7ckVgrwZB1FZHZz/wOS45WocFV/xafTGfTI++2nXDCu+FeSFuGCeFie9Lp9o
Le6cFmHpjW2CmMT2aD3OmiQFZjTJjyzT3PRZNGcIU23y3jdKclAaakWmZhtPTF6TysejPcxAFqH+
BVvydPHp3MIYxwnKR9GWiHxTZjR0aWTQXxuQ3YqqNNVcAYmpatKj10XhCKVDuDNPiljpQN53dO5O
ZVqUaHc7/guXTYojWlQYE8G/ZmkUXE+0SpiOTrB3AN8H4GBDSiHH8W8QtLyg9u2jhiJsxaKEo5pK
ECjKEMb/5zEzRt48psuTFRm3qYwYz+g48YT15NdYzb/9W8iAoslfN41VKeb2vNK+8sFOn0RbhlBC
F4k5yEYt9y+nGdJqFhnfyiwE/Wk354fIGddXZ0n0M0OhBPrFpIqcq+8bzLpLEA/Xrhvjmrw2MiBO
C36e+cV2WdcFBisDjpRkfWjuo2Ki0l8F4fT2CbBiR/XF2j3bIeoyOv15g3BqpZ/dNSNS8DJNzEzt
aMj9aho6aBCnlyjZ3X+rJTOLujHunYXVaBjrm2gfPyFZKo1gZ0IEKmsXa/WwVw2hJeGOSpSiod95
zqB4SDDagSmHn0/20XVOubXgMEwYy4ZCuezCPZdwy6MMD2s5b7IzEBqxXKMD6ejBhLl+wG8dhBZs
wq5bwTcTUNHQ07YIGnEihwcJGTQIdq6NSL3cO3d5CWG1npATpl+FW/dfL5r5DlunbMEfGKxfjPbe
MRtbVZzMxa/Akx4aRfCuHptCXKOjO/DVCNpS7Dlq7gzGzmf/ow5EeQuVtsGUwVdbyvxUUqGYXYj0
86ergPzkRnHE59FBB3PT7HJqk/VvzyjTvYEYyTJqQv9BPnD1Lsd0LhNRRxAlVofAjbgYNNEl4q10
a4jiE1SlOzukcKvQYhVHzDJoAd9+CC0JfVwIyC1Nh1g6CejZfT7rRWDKhFR1JwxyiVuqdMAQ0tb6
Uj64kKov4J3zUOPlaZyydGqFECaBv4cnz1kENy4jVmy9E3LVWLJj8Nq1B8dSJN8rpkNFczf144Oh
o0lrRplPvtUrxMd7450HBRXVHzqU2j0ZZemNgWKaoysaBiaXsX2t85NwcozHkS4uVPdxXWPTl9+U
vcrn86cpnaUi4QTG2yW911YPORy5aIUtZVHoKAgfh+Y04LMR0st3X4xSSCcnExyvCc+IXspVDSI/
k6yojwAnCYZLc6hSkqeUSIh5D314N2ijtOUs59Vhz0n0HSxbzoGkhaWncVbxnU+ABhsBx7j1h5wt
DgCsRNtHM7gUtM7Bbh8n4smCztODB/yeQ7XTtvZ8fNCWs5g57hrUFHFvJRMVpJQOS4nOZTj8euUa
MGglJjEQk2S98pkcCEICN5HC0rPySjigsoXI6JAhtYY8sZylga/x9IS/RujfJAF7ewesKWq50/Fj
ekEprZFH4e3lQ9VQvWoFOgaf98NAvSLennIqEi/GcsoSl5NBSUMtaUjK0NxDDJJYk+7DT2Ezr81v
9yXscYIfYEp2qam0rqGc+HdKa3VeHN+/rQfhNmwCDIM/gvl1Zwuk6JCbFMBWL/AlN++545NQ0I39
U0Ad937xjd02V9CuCM2iT9pOZea9DXuvO+40HKSRLTVS+RXqmgWKCNdN5MQYsqUSJPZVXZVqh56o
sAbr2VH8LZmgZ5C2D2yj6pT6nbN62yQ0XpKt+Vq/eD5P2hbcuLxcqagpLfGl3I/cEuIIdFoyIDxx
QWQBUKQ9zbypcgXZcoAaGkuZgpaMH7CQ0YfgRizCLFshEC8YomZ2tXJiFMI2r0LzvzQUzS2ziXon
+Q3tHH5yk8VDLwr3/RxeJ0L5Rn5E+4GhBaA7ifZ/AGPWcKpACpNCaQgtK2fUIg17ofkFeQwYcYu9
8BSFHtFjBg07a8IzABnY5koTD5/jzB9XZp06hyDQJUy70GzWt+WqUXKejYfvvq/2AIaqD9BaymgW
1jmlbW7iPT3MGuPmUuBZPomO/qUv0f/i+baq4H3qz9MZiU40eqyTEmH8D8BEPlpNLjE8c/MzOsGO
t1OianZiqQLf+bwgX2vAYo2a2tXyzOijdqJJE0mMCT0htK51nG5tqoOj7TNq2cczEp/Jsbdp92io
dpLQKODyxD3dLim0oeJiXYfuURe5QSlL92giv5Wymvin+m3l9XoVIekxacNl9DKVzG5oMKfeyz8A
iATeV+YI8TYnybl/VzA3CIsn5qbxUt5T73HP8A0Ka6R6PxAP0lZfUZlK6MJtt5Wz9aZLWMXcTcdw
MbxFBLsuMJeFJiM1+QkO5BcV0zHjn7yFmEkO6A9aqNl01DIvbZ2EAeQh0AgWUzFPaI5RURQHW/6W
dMq26c3z6ondQs+rP4YFzYbjncv6oD82RBRwHbG0tylZrXnngimv7kIolowL49pe64Dy360C8txE
U3/cyaLXthyyWCaCaDRfln7KE2+LTVbaNIyx+ZH4xCCKJMAoePVehBlyPohiLw7zJHGdGzMOYYxY
FbbkQJhJLZ0KYw/10V+B2MLxnsHDJG+gueGiiisJCUAT4bm/QyEvnR0TI3O2Le5moW6auL84/KS1
a9MpuaIgNgmuca+B0l1ZCaZXLQTrAceftIlKbdzB6Mb8AQhx4jocZLVoe5REVIskRaXna4UCaaix
SInut0SzL3FzNejLMaRCCAgkRMzitHRAAF7i/uDlX4Yfb6UEv996g/keYnB7GsUSGDLwJ8wuQKO8
BlfRRbPnnUS/st1a3hVSYeAasUs7p8Tv/rAitb5HgDyfAztiTkC+g18LUo2v+VEN7x8GvrZrRJMX
iVocBijb0EUcQWdMDVcYKTlQZHWTkvV1JkgTdbCb/PTJs5PYZwb54FU4uzLIUUGxRh5Afh0gwvWu
DX5XWtrqNudPGQz6hRz/KOvdnQQnDw4PFYK5cvLMuI0xeGL9DPp7ues/0XJbLlWwYD7JLzlac+Mi
KM4GN2JJz/s30MkAddYHd/gEKS1FPrLYftGMLchrvw6My1jeIPSxpnbTC1n12KNLolxO5oNj0lRf
1Zk8t7xvKvgLpIimF8zRVWVslT4cooUpX8GpKfZuh4pedeWAiO7zvafJh4cU5NOTcQ+ebHVf3qf5
a0k4VMAleEf0TtP5
`pragma protect end_protected
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="default"
`pragma protect author_info="default"
`pragma protect encrypt_agent="Synplify encryptP1735.pl"
`pragma protect encrypt_agent_info="Synplify encryptP1735.pl Version 1.1"

`pragma protect encoding=(enctype="base64", line_length=76, bytes=256)
`pragma protect key_keyowner="Synplicity"
`pragma protect key_keyname="SYNP05_001"
`pragma protect key_method="rsa"
`pragma protect key_block
ga7z3iGMhGhga7TzPGleypVOHJn9S7KEP16RJ6j/y4QGRddc7/SJdXJ2zPvm8FTCqWlJhu6/s34X
gPP3kw7dN1YdiZ3wZ0Vzt8uhC/B62KTkMGylsJT3Hm/4AVsby+VuOus10FHgOgp78G6FqJDW2hD4
FEF7AvpJ8kF9S1ZR/yBaB9R5/vEzgMTG6H0b1hzTpBGPyaW1S33KG60mDs4uY1wSc9WkIOuDsX13
gE5v3E3AdV0s35W8mk90srPFan8A4v9WhQvKv0pRdTPwajKYNoHYw9l0a0ijfdCCo0SwbSJr+KOr
7KJQNnQdeGn2Y8dg3BGFPO1H0k02bZuSqUQ8rQ==

`pragma protect encoding=(enctype="base64", line_length=76, bytes=256)
`pragma protect key_keyowner="GoWin"
`pragma protect key_keyname="GoWin2016"
`pragma protect key_method="rsa"
`pragma protect key_block
dBwrqXpaPIvc4b2fzIcAYNKycDBKm/hw0N9OirP+O5J0w47WHpIJLrz+YZdtlXZ+W2OT1CCdKga8
l9q6LpHNXfMJe0tSBaUQJS9kx12QCBYd7pz6Zz4XteULmwejqAW/r/1SNtjKdsFfgoOhPbvsYv0n
RR9WE79+rnvNSo03sWloLz3If8EsTQUj+4AuHA6W5eeLCFFrjEJDELred9ftNf+GjbKQ4DD9VT1l
GYpqKI157tMW7VzaYctB1tIYsZm6N1scQY5/pen6aJE9XG/GVJc/lUhiKfjKkAB4R0V1b6xO6o/L
Z0CvpttfY2ekIVc0VuCKq5gMTfn8BkW7RjZNRA==

`pragma protect data_keyowner="default-ip-vendor"
`pragma protect data_keyname="default-ip-key"
`pragma protect data_method="aes128-cbc"
`pragma protect encoding=(enctype="base64", line_length=76, bytes=9072)
`pragma protect data_block
3MLlIGXYAu+SNVZUrN9axPWxB76fSavWP25CyQigoZQ3T579rH2tX4mOroKAFnY6MCrE4zy5SoFT
o9pFhWobhy1JNncmCcy/a0fRL9ZlIyjwjHAt323ZL0R5G1zw5cvTmFWPoZX0yo775l85Oj07XBYY
i+0FcCRCKdgsQGwhMUnpc6ET4ttBmjQUuxB6g1Afy5ISJRNYs77D5E8aOFrmzUzDFsE9BGcX8wUT
bT4zFmjkBZBQ+KrbdhaUiVbninMVuzKJe0egFOCGcc6CdMPwZP2SxWGkscRsjPCAUdXGIydg5Z31
50m/zUoKITRK4jViYvnHt4f6sELIUTWEwPvxSg4M+j+wpDH8hMQC98bpm495w9Lz7AbFBmLBe5IG
17+sbfU7k0MY2fUrDvsniZvkyXNkbKvNrkm2E9MAmf3uKtqsnMU/tF2um9tYyMuoXrnv+cf1WHME
rcGa/NDEnGr3zL8P+jWgeThli88TgswwgsRldtZSZHdEDO1R1Eb97kPR2KAaazYlo2Q2STr+5F6V
SY1q0ie4TtY/nmeVptSZJNGauW3hhgmAK4fuCh0LfgbkBsnHNuCX8t9sRAwVUkoEOlvg+hIeL3ch
IbMuCTBsi9ym1EZ2NwdIt6YMzhAa6xgt6mL0uQSzppyrK9CSimYyzPbah+kviBaNcZ+XJClYLFwg
Dt034rBFaffea3MI9/T6EckVHZwmBgwvpnfxe5dIdxVZcMCrn14d+8gHoeJtodrk7RCejHv+C9Jn
yRjIaiu6w3mbAeAL4r66PbCB+S92jMdnwdBtSBcwI+pRfl8Y1ZjnMUax1D4+e4G/2vS04zWOHJPK
TAm5M/l7TRLujzCl4M5tq+MN/Sl/TrmT6Z4/ZBXtoFpOHicvprtU+bB6bA/TDiQ+wyauUCUWMDnD
F2sWssLTcUSqWyGH8nZQJkJU1GRznsjpDp4OUZFEoGr1SIfqUXOeUdRWE7kTsTGtuLLkFRULD9ZC
icKwOzgQXLWvy1haIHsyX6SZ+d2z16A+qjc4h9yGuTAjU8NLa0V/nk/gnsMB1qd073hph6QLxLJK
r4sFXdYNYgCk5RaS44kcalofpqStJQULijgevhq0IIAiHku9ZgDSCzWAw3Mr5M2bNizLX2XXA2zw
yD5SKKgh8NLJ62Z1MJq1d/+XEurLezROXf2MzGpmtx5eT+YNTMToyw4wlcI7tOteLNTVwpN45tUQ
B+wyQRROLfJbya1slSCz3CBx0TkfIQfh2iiO78hl2uIlnw7hygM5cDhSSbRATA0xa7ahqhvOPN7M
cHlx2JtFdxdsqSaZD9QoJ639DDyU3Hou+ECwMn0csUSwgAS8rtGVdP0Of14CplgwrGPXstO6akKA
3u+imfQ/w8L/PLKXBmZ4JDbURy7k1H6RKbw37csxd/ZvrS/pSmIkcNCzp/c2DuOoQ7gmrvF/T6P6
o66nwV4BSbtkXVm1Gd6pj8kuzFas4d8qUgIJYtO74n7f/EHBC4KRyKr547xiGiwhk9b9qd0mjPKY
rhYsYy9gXuZh3r68RGneNEq01MvW6g9QFwK1ZOIvZDYOR4QWzSf3jaria7TfeR04B0hTDmN2pnIe
G0GNQyny7szBaDLk+3oC5dKi2x7IBMiFePNumBGpRQwF3BZOBafJAtsThr6J0+IuaIyGTu6q0CRE
pK6/stbZUIyDHLZTtsEiDvCUoqJt1Nwycg1jZabyqczbNym1H0NA+utNZBXESxVE+E0tL5xp64UF
6UUd+qxyLwKovERkzivDR8GuW1zTirEOV5S4VxepjAekJHQRl/DLLebsO05p1WmBlr64t8l3I2Z4
eBoTyoAckywhyY3Hef2UK2jwBO8dnRLD1Fu46o95g5M70RM/CdS1OdLKSF5ccJEDtzouHFkJV1Uj
jF3ui454vNAg2ROOQ3kKuyo5BsEY2EVCu3TpZq4c/q9GQLsRGPOnx3VcTR+6BZb9QBmDwr5qk+/F
Mfy0nKqqzp3OK73AWybRMjmJczTm6ffP4zxEkfUdzR127EO+OljvRItBn8LSuKgqUpIu2NxDCg+f
A8xmKgcdP5Vj8cz+tus1NipaLcnS3rd6rslS/DaabQM/fOpx4ERbftZUSiDhPxRfGlVjhYH1zMEk
pr486KmY6LfVGaqc2pCdgIkuSoohsNiPN8xmmK5O9HjxRm7IYdaUIvotow0YeYsJys+80/gJB5s6
cE/ss5YkBWNMAqtri10qAqP/lHRchjbTFTFInn1auRmyFcN5WTjU9MqXhbmBIpJrVs6hQ8bjrGbe
udyynSp5mkE0eE/e2v5I1wi1YhxlXU/wpSQkq7AW/DgOKirxvaKomORblPuNuqND5ETjQo+jpEPM
80/aOZIyPqN0aWmrTJE0jsjxS1AJ4MOENCzTG523Wq1bgye8XzrN4fo53VpdHD6EPKSh7ZgGV7sq
giQ8mzKHA5CetG2XXI6zrPk7Oe4z8m90oe+OF3HP34C4sTOp/x3Y+GqefIC7NoHPNtvs6PK4n21W
QJDfypWh5VF59VtNEgflzAT2wYDVtih7VEgDNBwrj5ychDhaeRx4+0dTJ9BZTa/Q0qZqOY4erpsq
jvneKxGNPh7zRngog7RWOBuH1Hi9ahuIiY+gEC8RxoTw0q9WCloHfF6cK42Bey41W7Nkg8Ic3W6O
AV81HlRcI218/r7yKU/7urKe8KAq0lmfWI0uIobow6NRr57vlBBhnMIl/DXynMAD0MicHsH1Dhyn
h+XWBoQuDUWkaHIh4zZ/+1qRMEs0NnSiSUJpOxoccGc+tyhoKIypXhHvUevk4IqtTmdXqAG9BJVV
k5OY9fhhlE2OW/ibdkZv1N8TAqzbACTxaJsG4yd9IXNrWQH3memdIJYipNklf5EjC/KvbTm5tyl+
BLxlplNCoR4T5q2klsjPNTl8nKAiMYCZJ29rISm9ghJjvtpxxC7iQxNuwy8DpjfL8Uf4MMBxii/H
GSJtEZy1R7DGqeOvCIAWAjS1+kkxdMrlh0x3ruEo2+mWagYuF7zcRwv3TrcxsdpZpxjAK3KuJQ5d
X94lkof9p94Q9FjBqgLyhEjFTPbeSIdMHrEiuPoqCq/SHstw6UAe/HyD6+3m2O2WR1U2m9uPatvm
sJxRvmVVaHWurvpn1JNRY5/mpZqXlkjzuf/rk4eL7YaveH1F0WX+Ql3Pd0MA4RpPOCPoYJ6ooi3X
oVoBCaBgNLwuE9nJoaTWldtbdFa4ZaDZk7rQMlAKVWXu5XPEChTjxfzXr9iZw8Qdf1rTNBPLxMWO
LS48BLsmr5GXjy67UEUXHgGbVRrUX2AYtWS9hX1O9CEOcvgQiFyWG7+HS9TBB6SQ2461BLLzDSIm
tHQ82QNlJVtLqGTo0WcNrWtZBNk8qWHaU3vXA5QOlhzZmHw9E/y6jLn511lV/OUgJnhM+VkJUv5u
1GWSh+SGQ7IGzBlp1mAMXXSKsY9cSzVqiU7ytCkCfz7j3DJH5ntdAicnI7krHr+QdHoHVl3cPRNN
NTik7Oj2TIhkPWTVsDBGPqiRUwIeX6/EI9jZpwpEEOFrirGLMXLQlE4bDVag+ARha7L0G1Qn/UwS
ejMGqfZQRAgKydtDRMPe5ZVBcXjxlbFRxDPhda1EEu9YwjoxssFUFYaTKNMkzgd/ILMYuoWISXaK
+L64nS9GUjgI6nDexUaG+DxiNSa9V3et6jDkOQxxrgWcmQBpkk37KtycdmM0jrStFP5wmOsnlJFp
SCGPeuT7Jqp7MdnYaR5o3vKVglmGTbwjVEyEhlWMC2Bbyue7NnT/dyA0LgjQbOF69e2BR2bdmIIP
aBoT0VEoRqavKJW4VVJaM54H1gcMOvTiiwzgnJDFqLa7/UA/7wMiCGu4uBnB3/kQzacm2hlKuJQf
T0+vWNMiVBUy2cr3ft0/kuEG36VBq+hWxfKK49u9O1qhxvIIn1z1ZWZZD3MHuAZXojeGQbtv3kru
U3XT+pJVLh5oW7JXXxSWdaz2//oEhs7UgNjE6GxBsIMlGPBbkJ/ycx5yfyxee/gm59BlN6y3qJxe
INbnePJ8joraeLI54HYhmuIWx90XFHYoDJPGQspHtIFbLkbuwDmzVGbD7LA5GRjFnNUrTZfAP1EV
adRX/fDuSPpw1emPPqmQZH5VK30d64GZveWzK9i1yfrdv5e65TEzX6LlxttTYQKkEP+dtczwig//
R1YueNMWN0TwjToe2drBo7oIH3dvjjmCJGzj7L0KVXsa9T9OWhDmY3bFcKwLDrLfrOm4R/IuFEHK
WOdLDSei1hDzy7wy/K8jki8xgNIqCnChyI0UL0h7MGpoJZmBKzpmB21NrbYCdS+XnclyZ4pPkj97
Ylxo6BmW16US+sj65NAvt7uBNJHj+3T8wr3qBqSrSQsvZLNHSB5/u+5ZrPQSNqbhhjQv0NxUm8rW
8mlir3nvxXFJPZ3K+S6GI2Qwnf2OY2Rw6oMPtCsWx/sQiTfPQtb0pb9mnbOcVNeiEbHXgFZ0MLGz
HSxuKW1kexbxYUG3eu6vL1dlUHRKIQ/2irLYTwymVewOAwSODl+75/uB8Wo0kVVvpXGw/mTINAYu
7qVxHRYXpj/ksW4pfMUjP/9kM80OPdcSc/1g9yUPA2RX7QkGwH4JCwwFsIgv1mvu601jFz0O9Bkl
0PpkocFdGAcJZC9DhmjGWZD2cCN9j8QnvkQzeLUERyt2rqFfavwGkaLpxkfrv6OpLM+hpop9o/W7
f/p/JrT5qiANXTGmqz3ylmPoU7Tu4TIZURP/95dqi3BHf6QvnUPTKGAl4uafN0PLzeEkjspNN5/C
vni04/K/QKDpgxa85gtsasDqyIKmwUwKZM9db8gdA4mIUc8FLdgw9dfgKKI4tgB5EpPMO/Tj4lis
tqjm7rIoMX1dCl02nm+cc00Ed2SnpCSRajJwqkmgz9Uw6BQK5BquKLHcV+uKhZLq96f6F7NxXbnC
VSmpjLjMAEWoUhzZfYGWzNZOcaJaQoYR9IXGrPsoNr30J2p3o8wNrqGikw9KYNxK2WvLCY9Mm7xZ
ANoDsp+v7SBkr8eLvaW46it+Y7rYG5klsRcSUw2nGHzcpwmn6qcJp532CjFhZ8hmxQdCEJZIwILp
uVzRdxU2t90fe9mLoXkrhCopSuvSplsAbKZ6yaOhsSOu4PuU5VUVh/u6OF/PfBHMdXgwxU8FGb0y
hUR83gXciXE6dREXeQKuXfCaGYRt3sEnSdXhFFTMqzCvmb7EX97OWDNl2ogFkF1eh8vEFp0cO/9x
ayCzUdCED5U4SZwamqb/MDo9zUz0PLFfyfocYTFS3vlN2VJ3g9+6zxksTm1dsSso6oHVH8ZJP6wd
KIr9m8QKTd0FXZnWiH8hJg6E73Ssrjj1b7gwI40w3m+jM0O4LqBgHZctjoM+4eYsfe85yhVIUyKV
Urgl0O4NuR1uZsW1VMGVtyngNkI31gbHIWv572fxN4ikoANmSxhGNAG8/qCWyXdQfJUNELlRqqQa
kAwhWwDVJZ+k50DJZTz8jARz55BNIjVR8ErTF/GuvisBZVjiueUM3GW1QUQeP/jr86MB0LIYNccP
7DHwyT47vp2fhU7IuvD8FiP6/DegR7eAvpv3T+B+xcT/I0uB2x8fDgPJw1/b7F5HfvZCIbNb5SVH
Tw7kBYyOuTrwFrANCDbsV1429WaRXUdBnqS4UbNEGIFXNSPuHpR13Ge402Mxb5MyuIoWP6pRx+Eg
Pj+pw3+oMLd+I+j8zxN+qdK0FuoI6nIHh8NDD61SHNGXSOeWuJ2wEGqziBE6o/rm7lnw/bQdqxSR
YV5Byzql8lSKdW32uiMMYz5nKDMtqxStIVSJkUCxjUlJ0mnGjcnXo5P7leZKY58LPiS94oXhcC1O
kzKxrKVJznqpGM6Eln8v0BX2ilCKY/b4oLhLU3B0u+qFUU2olYnVfQhZM3E1Tp5gS54P2pdf1v7c
KMuRwNntpy+X5hZYMgazx7Dov2KLO0FXoYNaiIj/o15wKmxexJw2MwilFA9cGzvh4CMHx38XNzKc
wbmBHeWpHQ2ARcOylDwPaiSrZ5E5d47fg7raWfP4ysjybfrEWn85I6dCXk6w0qhPvAXOiW4AZ3bh
xgXiJsP7o766J5nn7rYPh42eWEfuBRnR8dh4lgEAHrSM0gB69R5KiLHVQ5/R4XG1QSCw4SsV5Wuo
ths/6EB8J3AY3AfdjIkHCCeVbt5x8c4K68sXKhTR+ifR5K+G5ToxIAY+OhoJ54flErjCOsmF/Wiu
rfX2Wa8sXm4npR8kPiC5at4zYcE4qRzc0xiEcXBo9v8uBV1Vifu6gh4z5HlYIFA5dGnrDkzIlSIK
dYpVB9FND7PXET8E0tDhT3Flaubox2Hq5oXdATN8WCNhrjM4V/hELCobdz326sZQhR5GUkDcApny
8Tu4F2YAlvhn2A8Ni4Rj3USuxSiyNiEg1PAK3+1XmtcJjKSIl4wJRNu3+Jr2xP+LlOpkl124rb6J
Je/Gg5bnxJndk1c/DuCX3w7v8cZrwLv1uAZ/6bzHmHGswjZVzzR1xNmjDtRzChlCNkuAEz2kRbLx
TGi4H0rYWZ6AR8ZksqJiY4ufxrQg6Ldr8WBUJmMvtPmytfptUDr2j2sHyxEQFfzzya/rhjL11VKL
N7QNG5cVC5N31XO+mpdD6mn8gvddDzOl/qRc6SuOJsMjfPTbzBexpAWrLA9YSaGy/2R7d9hDZvWH
f5qEB1TRWgjyyKuu3LEVeIMTJgnHmeCOujSjgPByFLXLpFVmjFDrB5Aq8cu3WtWI/NfA7Qem5gy2
xsEwm5qpaMi/nT+K4rQPJ1N4gMikPiIoIGI1I9NSxhJrh3PeUJNOh4qrXWU1Wu/XMKwZnPCe9pak
HvHKNuIrD/jHS7WIas9/1iLRBIonDsenldC2bBC28pf5z3WzOe0WPpYYaGQ827RaH73ls9i955f7
qkA82W14/tV1nEVK5kYtL2JaPDbUU6Mfq7liEafhvOXdTnHAKAykh9k7HNAniy5DUH0nnOe3lVjG
yr29Ha3farSkRstToaPVDiM+kHJ8N+TCwK72uI7LbeS2+2LQRlVmYo4X8PY/ASciygc1olGkqFh/
qMNFN6cO7zZhDXiCSeSPwyvjeZXiiGBoH4a2w8IBU2AX7tG5MDMkudV+spTesytgJcAiQs6CpfwF
XsaGajW8R6h291d3smw/AY5JVSjZsYTSvsjofb2Zxm5nd5iL3iWJXoeWWi+3mZQGkXW2BMHF2CVS
71igJE+ptLEY45GJad81yapgU4axkimT3BMSoPqNfhxO5OV3Ta3odZgdYhdqnP+teV2RG/M2Hd/H
E288O8tfTHu90FcsNy/SgvOzLmoPcd0/jHLd56BDI4zowvJ69W1PZyNi2AgFDDHSY64wVDAD0Cnc
6nomSA019TnER/cjplfR/my3/bQV5gcWPTh84/J5wculwphZJOuhElTGmOEhV1jeyaq1Fd1hzTTs
lDb6D1sOMQmeA+lhr8nVt4CThr6LEBDzR0DwrW6HQCfElBCaWqCbnWiKiR4gJSIGEzIn1YHKLcCu
LfEe57KAA1/tUdDDJawHF9BsHlIPOdLTLTORxyTMSOspPtX9NVSGGUWnVvU8FmTNgyVplcWAXUIT
ee9Yg1GI27KLGOkDIezcY4sXmfonRF7zo82INxyaGwCGcRsv8J0VnEuBiejsOBoyo/8OrBH107B+
4mAc3+SyCipuEv1GGPGUbQSbUFhd8bAFZSgTVO223XsnTnv5ewREPpjR9QrBsdWdEKtHRSxfwqbM
mtPlrN3vUor4eQP8Db4NpsWWkzKRD0rVDSpXhpK9d7HGXIHpk4SXGSM9nTh2+e8N/SFKI9vr5mx8
NwwnSy4d0+wgkNtmxRUXUa3IiPFHU/+hE3CDn/4ntwb2GlKBRD6Ae6Y1ehUydDMTz38WN6cs7mwv
juVogt75j5Nk8CmgaQMwbkVFALve36moW/zZokz4L7mitltlw0/FYgtIAe3hqBryx2rQvWDf0C2W
Oh4lru29HTO/+aYwUubowRlHDa0/8At1XdjjdkOuy8rdPtGqpI0CZAJ7/DqNlAPa0gSfKT5Au7kP
YjYpg+Od05YDKTRHtEL8KTagsyy1mcf6P7W+75CEdG4k99e3J2UIXN59F75xz37cnfNt2zwWo8zU
slA09I2lTSE/zMRFXLwpUL2OZTCm8sTOfJaF59d767021lvzPdEnJkGrV2e0U4rQht4rm6Nx7NfE
Ki7tT5Rhe7FyvdRAxRhjmY1/2771QDsWk5mnuOrc4cZz63aJ/cxz1d4UJNa7TDqO2Zinpr3SbAyb
6HYsI3502PxmvK5mWOxRhmbtA5dcuDOFHSCvJkJn1Fim185yR3CbSqJ9mnavtlCY+W+hHZSUVg8P
syLhpJ0i/j2nTpJ39m3cYrFYGqRiBRf3ZDHOn3VFxfWqXpo8WCpeh2cm2yAL6Q6FBMulgN5Z9gAt
oEvw9gP+CTbAiLK4q84JfvUWssnxx49+USxDBjb0IlqWNFGpzv/JQE1jhgELytU0IsPHKFXXug8G
TXYg8h/HyNAKbpnhDyWmCJTS3Z5AfwHCFT2u0sAhLQaeDVFw2DU+IHWOcnkSfnbHElFir4Hfu7rd
EwOcYOgMs5rDiaiTrZwFkK3CKX/1kyMs3S9IgPKgrsXz4uIHvTMzZ3hQYXTC5Y4H9cvlN2Ax/ZRC
0W85mvpe26738kQ52yzmvf7eqJlgl1cNSNii+RWbbZPbk3VhTri/nlMmnwYMbD5gjWBY33A5gqfO
sBDn+F2O6Q6rk4M5WBHKAFleJJdf5IKSkd59TUsiDZvr1UFZCv9Ppxt9L6ZMPy9644PmqeX5TVzT
YeOGylwSDlWtAImiUHOWL3hxFR3XPBou7REWQHnXkRURf+MCBbhOauPVdHfwNkry3/ByP5JBD3RO
0BbSaWAc1Duqhmfy6me5oniY/6iQg/rrtyJ3ZG3U3qLgExk7tn+qxHRVV7sb84TCUojRsjdo+DSN
gk0uEfGVS320FuP78CH98RhDObVqWkjsjb8HxVbFShRf0wHoXjGIYPvSnKrT9VhN+VQkKCmUF7vP
48eq2mtrbmbOlfdkVMSDgUjuMHKhpN7/X3gKEQRaB8ai+luUtEXTKgF6vvt82XMOTswnQmanMgha
0ENrZ28dHSwgE0Snob5mYlafk1QsBazL9KuWopmgb4WsXVR9HxAkysmOa6QShVfpMXgF/lurt2eK
7zG9GMPp+451cr6BwWxmWtN9F30ZuNN26EV6onk+WCuwniVYsXJu5GJl2eATWA7gT6yNcwlnAW3V
N6qJ5Ce802YxQyYHGqr/Dv9TRswto7rNGkIkpVTE1D4mO7zyr4Vby1s/0806/bme07JVbOUotqbC
SVbJ0/W9m8tcKHd8jguDPJ3Wo2Irur819WuhbS9i1LjzNjsckztEWJKcRuCslVYfcrM8VIH/r43M
WxzbhyP+bCshRy7wEImhKIWowgsqM2NUPjzM5GY9NkDtf36bZmYZjvqyA4iXuAy+I5eQKVykV3GV
nd8rbTqJMumcSCIoB8T4EiRkEdX5b9xSrpBVOHyMv+LYnk59mP+7w8WSeDfjkIGuUPpg115vexWa
3mP3L8c/qh/AAL+/IT48uiO8fyheRJ2IXCSQwe1KgTibe6qeCPLnPWg9OutX7ZOENh3f3C9HOPwc
G/Vdf546gc0Ao4Xg9HiXlbk68HCRbcV8SrazEXi3nomQsiTxjv3ZDOQT3yZREypy3t2lJp39xG5e
x9kMEc5NSczN3Sy11zER1sNG4HxEdMYATQaYUaVp7gctY7aRUFeQLWoWulNSVvS7+GZOeHMkHw5/
yRlZwGc+cbBTXZpE+k88139MNA8KTFjmInQ/pSK4gRsUKnOSChFGfMyVoxV3Z3603dBO+eTDGCIg
sqkfNZAlKZy4ewZ3IDFw1R0HQfctegwFKqK5k+b7qfP8TbB9CPlk2XYNoaQ4PV6fKlUOZY6lDZYZ
DaNuEsxmvI792YipnSqZ+NyjfOyyCpH5DXj09Ol1XKNESmxOzpsXSaHKJxV6Dz50wZl78nfMA4WV
uJnsePvE1g/OGZaDFZX7pPEFBcHzHoQ7wa/lPUlxhTuDYaCkytVl19ZJb74X4yCD5SCY7eLuOZ5J
f0zj7uwPjnLMu402QSr7htXY78j0+MhoC7zi5vUVBeqeXvw7vmsp0zxaghJ+DGJEFei2+ROSKqSy
yWvn3lU+b2GvYmpnTWY6XB2MAHuAriIgJ4ruPQM7vf9Xvmc/GolxsRVr/t6UH4tl+67q5X+Qsr5e
eLBG4eWagKTrZYhLeeIhbsYG1ZuiOGJYVIub4e+StYBVEGtCfLzB/fJAsRESKF982kcbeg0M83t8
3UYhH3o3OE2vQX9ez+NRvo5IQF+wivGT0SK55QeQd/fRktmwSBHxIiB1hQiWy+GPj7hwHJs/SROW
8Ul042DLYuUKLkfgKNnWp6A2QkPGvgTaZI5mD4sU6okw8hErv3KCMrtT/DTepa0vSCzaZkfz1D0n
0/6wdQ0UNam4BKxH2AC8FPyVcbOdzlZNiNLUGjDMMIqoqDAJqK0y4gykOMgBn80S97VestIWSCsn
AFFReSu4bCLu3XlH40qljY6wbCw82dEgX8zInQ285Xyr9H9BnpfC0yYVkuNTu5a8qFNVEpc2FW5N
1xHep8yYN3nWEpc2EKdOzDiKYpOzXlsmrqDY4lgGiQHKvHzYSMzlBUgQzrr/eaKeeBcg7lTkXIS0
uE9xM1Dnxrjz4/NooqxChQyRsqNGIxGnTDEZkkNesW5drt32z6ILExYiTPVzNAMKMkWPxLrz5OZO
/RDWzzMteLKyzGbRrbL0UTJqJ7KzUIFO287TnxLWQhnmk50OZ1mk/ZPWebYjtORDeQ/ksyoAcsT9
FOeAx0Wg/WUpMjUC5rlx+9nQYQ2rVVQ3tPe9GnH/AGm/SFUDvpWQ8MYFua67HgTCbEzWJM9796Yg
xff1U8MwYyGKMajYwTqJCx0LvDlAZtH/s4Bjab0Gb/aRN1kF4mE3tO24yRC0DtRyGX9DV7sx9T5b
5EghNagRvM0iftiYTaeJDEKZ95sx4pV1/ITAzm1qeoZad1ybAiiGeqmAzgDuciavuVP7TtuMYiGj
DqxdbI1ay1UVo/e4DfY1Y4+uu/EtFj9DLXKD1jeEtkYPgzgKIW66JJarx/6BLgZX6ES5CkvhU7ja
B3FWagRY5+/iYjRPL/R47vQq/g33VIn6pTp78y6Ez/uUv+LDfGe1J6TuSdZuvhNgyeU15VnRKIym
Lhnm3qtqfv/angAozu26sbPXYzWb38h4dvZGwUZVD/a23013aRTClLJy+QDiRaxeGgF9bnXh8jfg
RnCAYeW0qRvv2DgVRWKFjUGkJQqRfO+wMd+s+iY38Us+wcTD4qWcdW+SgY+7gvA9R60FA9g2Z1MF
c0XSHj2NKu5vr9ztETZjqGJ46nkpduHBoPL95u7CaHDfeASF6yoWxgLbDswJkfLuPAl96TfeSMFL
8VG+f0VSV1EN/CL92AQqm0n6KczWCu/SLY/8PmY5sOTJMVz0dvRyV+gZBbRSPtixs6eklHCOMSzz
pekeY9VydYZEqQ11cmKULGF5/zNgA51lHjU6rRWOoxTRtveEyLiPz9F9zOfSJElhHH6b1R+MNkX4
WnLs82rY/3I/rY1nTNvTZcvmqGURL1GdHLE/c2WwSmWysp6hoitzNoi9stuE+6IXnuDahIvI/Paj
AjxhUbZ5TxlFZ6RTbaAaE8wn7jrp8wlBb9KVfw8SliiEYExYhdbC7X3zIr4+pR7ZDfxA/sbWx2qg
IjSSJkCcjuhnvzdLHBaQJrN1HmNUHYSQUBL6eolvzAzISiAdRNbDdJEtrYD5xUysTi1SMvSylURB
gWywb9XtPlZMnqMPDgNLpS8iL5zbB/mHbQ8HnYPXgHd2d8ecCLMKVuyR3wrU+sheD6NsAM9E1uL+
w86Z2P1C/UZygh3aAzBFK9/UHMAzM5K1LXxk+Gebn4AyFohrdVamFp/cljywjlrpVqFC+e864pGs
fuC1ghoEq7pMFhUOiiLDLI7tmw91bX51OD9hnarCl2zJmpjwLQ4dIKkexZFNTilP7hI7dw3HxvpS
CmVns1GH6E+t
`pragma protect end_protected
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="default"
`pragma protect author_info="default"
`pragma protect encrypt_agent="Synplify encryptP1735.pl"
`pragma protect encrypt_agent_info="Synplify encryptP1735.pl Version 1.1"

`pragma protect encoding=(enctype="base64", line_length=76, bytes=256)
`pragma protect key_keyowner="Synplicity"
`pragma protect key_keyname="SYNP05_001"
`pragma protect key_method="rsa"
`pragma protect key_block
FF92Y2BScS1tYCbOJ6nl/yrS9tO5nLdkcinIUmduQUlX/rEFHoa3Ivyk0aB+kXloe21LQE4kGkQ6
Q9+cOvbtZsLXojH8eCz5LSxZZmj1OY0HgImQvBdW/AXKvPSh/8qp2AkQS6z06aDmakr4JM27sgw4
e8FcV4tuRcqkGs7bb5nTeggXj+gCM8w1pZjupaF2huj2/7utBwg2caonPL9QnFqNhJnw1y8cEijm
U2tA1t1pCHmc/cfMmTL1KVw5knK/j+GUCQdryhHqwEoaWgcU/WsJ66DlhJyiBG8LqQzPrvznCBbb
LaJ3ZRAbBz91jljSVrMpulWLCnotPmY5QRPBNQ==

`pragma protect encoding=(enctype="base64", line_length=76, bytes=256)
`pragma protect key_keyowner="GoWin"
`pragma protect key_keyname="GoWin2016"
`pragma protect key_method="rsa"
`pragma protect key_block
cqAgpvQThUsKP1YQSQ4a4I/shkrWufEhsDBDReUcDIwQgy0J3zK8Xf8BMFoFrewCsS2KNDRzQ+ER
jCDGccgdbKH/8jqChdozG61idZWa0ns7506SogoQlXjlqxzJaYEQMyNxDX7Ycmqi2PkN9cXJyFzV
5txS0QofbL3mzPtdA044rsuP1fkQj0yHft0ysK4zktjTKWnJPMDoc1p9qdrOCvbt1ZBLB18dsflT
y4tm2j7ie4QPZbNefa8AuI4j7gxnCkSCkqJB+CSn4ks4ndlDn/a3c79q59d4UozEclqodJLD4obY
Qe0wLjtJvGaBIVSj8HG9RNO8kRI3GFa3bHt0Iw==

`pragma protect data_keyowner="default-ip-vendor"
`pragma protect data_keyname="default-ip-key"
`pragma protect data_method="aes128-cbc"
`pragma protect encoding=(enctype="base64", line_length=76, bytes=34448)
`pragma protect data_block
GMWtVErQpQVB3QwSqSu3WLxWBruia83TiqFim1P5yonkOBqD0gjMvU2G7mVGBBaenbnn+fnYB+PH
jvWo0y+KfEKZgc5j7VYN+0RMmwbU9TIha7v5/wTNogAJb6KmlLtSYphmoF8wNRarTaCy5b2nEHI6
kKTj9oOOPYDJJHgP11/9xZIl7g877hCKnUjGHY72ptPHCmGDuH06ny3wOp29cvOKHHnza45Qmsb7
1Z2nx1zIRx6Xy3Ow5FjzGOu6F+EW48n+NV7QkA96O4IU6DTe9hTU1IOWCTt7jQHPPLnS0y2fZvXx
7o1HwegqdHyN9JeOpG/RMLdmac7h9SP73Juxg0BbmNiSET6KwcnZYGfo3NNGBGIrLUtQLvm1Ak8Y
PVRbcVIjcxR1Jl6+IY+NruH+P31yhbUYFoVk5+dOkLzKf5wRlxGNVteAphomb69XGd30owusQK5h
zaKOzfxvks6nrdTchKhVMk0dKwLFeeMABLcA+o7gTMtKSxdZ803T9Y/GrrM3RciFK8Os6ci0CAYi
SIluySEYpDEUSWdINadQA7xSyMlc3LwJYfSZP6ET6CTGJLAn8F561cUXpjiOcp7oq6gpUbEo8xem
Rh6H+1jQrI7XIMLJ/JWUGOm1heyXad0gT0gwH+dbbZJMZkiHRPyEhcQI5KSD6DVeEjNQIiPPlazw
xKd3C9XNBKZCt/HhEy60hMHpi7BsbAwGSAL3fDZsJwU2OCHkIhFI5E6PsGgRNPULQtkHys+SjtR3
wSCanOV7zx8ADQjXGLAZgvhTUWGupHSSV6HbrEEPiUzSg+vV8sN7qGe17JvDcyRN6ADcu4PYvmyL
aH3bbCFHS86DtvtPM5OtXWtnhGZO/wZ8tqrbuCsyI7u7C9omHx3+weFTS0Ok/u0kv+OGiNSV/B7P
81r13bINRBBz0dT743FShzr7aDBAv16M1oOSBqjEaSKR2151mzOcLU18wpjGsgy76HF1fk52wLQA
QT+mhrCMPdvMIPaK8Z1rcIWr7q9a1Su4SR1BqJUNzq8/Qm8sCj2XsoKc+e8oUJ4ITPCHuo1BzQrQ
Nq12+g+WBGxzpS8UZrUZQIWnxERRXFbvawhl28hRURdPnKgC8/uXqjlC91rKesFsX4jMp31CNQQ9
aICs8mpFPQ82eBNRZIV00PoYJN601yVa2VH3jn9xELk+2y0NIPzSg+OEy3SPntcQkAl5CPjNjkHN
pe3Bv4vFSNGGS5Nn5qp2zQMZfvlk39ufnJBL02PI4N6e2wsZ+w6YJOseQq5nQP/noNeLzmXhKpZ5
9OSVHrZhm6iovRGTNjrE6YKn3FT3hdrzvicmsOBal3LJST0UP8YZ3bOri+MTRthkOolYtihcRsdO
grNtUp273INEdyMBmiLR2a3OAONXNfWgPUoBT6a34tWNELVhJ+SbQaApp4AnoNd10D3wYImMibfn
iHQBhbXsnYQNN3q84iSFjNLwXmnIjteXZjz3DDX7ECJwdWocdmuK3irOw5fyZErSItA8/FSvYf+G
xwigooZzTzbWABvpTExFP+wcfGT7zzP2zhGk4coN5IAI2WT9HIOKMez8D+PHGgQ8oNhCjwl08WSJ
5TdBkFHFKqm5Qn+5dmAkmoqCxgmZtoN0QffsicPyJcntbjTyEKjZ3KcXGxw9q1Jlh0Xz64mt/5yu
Mk6cFO4J/Mg6vO8n7/oHmukOdGLGXCcrtdfbwYQQWMpT7UFtjWLlrMmtmmLV8lXOask1NShNTqXN
FwBGg+Gq8yhNbckixSZBUrnFNfyIsDDGlsk4VRqMZbHvKAXQba9WTI4zFMtFYML+vBh/Eaul3tPA
8HLYmTlvQe+HokJ65NE9sVtYeXpmIsMqRTccyu6/loSs1FjVgsJcIP4N+cMWFdtWwSsAKb6F+C9d
GZosQhB7UC5HWcT0053GEa8WaNHHw0yG2zjtqsoZq+cZfUfV416fG//vLo5OBtofcxvso5+SbR5f
qrq7qL0hIVmaIbx7qoDSATLNj/5ujyq//sXLEhjoGAKxMjm0RSBFjXsx6tT2g5bCGD5ugLuBL5f2
1MKgJ02gpH9NkaH+MgXNfher2Kl7Cs971ZjgkHTeGFFq5TObpugWJWyL1aSZ89jmDrxZbBeEWiCW
4uf7lWk4mEt8aWYX5kd1uqdQr5TBK40z50pd8pspqBh5hqu+Ozo2PzwtYr+slMNJe5Iymdhm61ce
3Vkpj+qnCJNf3O6OvWnidumHcsB3IKYSosEI17qYXlOAc5K9g/cv48mmt27Frhs/UI3Np+cr6Os7
NgnP5M9QnSPOcc9gkxAPooKgYgDoysHHVDUef9K5q36jcZStx4m8xtf+rhuEwJlV3hEB80TbYcGf
n2nNOXLd+TdtQRaYhcROY4zB5155ljRHwmDGi00xNCWPKxyvbtMdVSDbnhhglANxHHFC9hsvEcSj
YBLW8trsKuI0r7LfGTRVgi01NfC/VmUzocMToGQWg10Omds6IXeCDZkNwK2d/p7E58CgpX8Orv3w
1trJb3EqLBpMyazHEGpLcWcsqWyy0K8FAonWctzV6730TN6ozaRVHXdfPrk1Wj7po1iU/V5Pb9et
WxTn6u7/UI8GG5N0IXovP0CviQ4fEVmfdfCtzi1o1d8hxW6teGPoZSGINDaPCIAbhnoLlCBWsbWu
tMEU3FIkXsCIzGM5BPYh04i+o+M55MtzpAGL9PmmbJgRpsS9Js23cyW1AQXsl1hOCrwASbJsbUIn
rzzTM4OcYwD4sttWzSsTIET2MbPfClnzZ2ktdrWdaL1Tp1lO8y+xftPXYnuMw2GGRDjGhCtKxxc/
eDuNHuLSO9K4a5IPaZlV1G9ndFhy9YfXiKWkPo91zpndK0AyGDu26IqK5UZzW5t21B9VspGjg3gD
G+/40OfHoHM9XJ9Oka3JyEk0QPutEKE9ls/ax1nGU2N3de2HVlRKjt7DwNuwFwGBFkIHb3sCenrp
RTyqbayilto7eZGAjTnSpBjkb0FIisBHWVVJ1UEZVC2DTo5So9CSqZtlZVaPmO/LviDOMzgHe+tp
5dWPP3DHzJ8CfgdSkZecgltfkhlSSxKsz9uCcHmDWcpa3r7+z4fpgGVBgVTsbTZomrwFdaF81Oyk
/egNA76akSyRqUIAe3BDJN1hKDKpGDo9b0OsUZCwh3snYJ/j/CrC7GG0mNJ35nVURJAYa7TTrPSY
XFGwa5xH4OiZLe6suWp/hlPv7B/Jm72Rr77Vn3Yf+faQWcoPB8kq1QWz4JgLBreLOOU/u/1NM0O9
dK/96CmsB0EY0lrY0VovZuD4QudQMApAagBVrm5tg1DxnUS9uIxy0ClBN2waif6NmuSSmtUhObQH
X7rKVFOvL9vicozqO1XiFh4uNmsxcOpR3PM2QfVS28oDAWRN8OPQ/N6HEq5jkjTAbBvOGiZD0REX
8h9r5sr684UxXrWL58Visv0kFk2X9bdpAEtxkTjPR8VUj+YatiN/AB42hPdKaR3yWrGi6MDl7PD4
8J1ThNee2X1YqbRR+rXMQx6etvOzTWYRmguGZxYF1/J6erAcHcAwuB9VOh+tBhUVXJgo6MuvPnje
blGlOI7Nkq0/SdmOdwmy9vwFMRcQoTyaKfwQbboOacCXbEtLC38P/p88yafYqW5qvd0njXA6zVGR
/ueu+NexbRS0XYMniwe23BetnoZ3Iz4Dh84IByo3BG7Th67rqnX0nmmyOSTgvoOcqyK1hIwsdrJq
ltYDewJ0gT3uunRAcyQQp4h2usTbkQTOwm2dj3ZEdqIuGlDMxPFK2+LWAdq3Qy/sVHGcEyDSegxB
mFI6g2KouLz/SfCa6mkF80WLOYi8YRnwNdl5BXCAjd3+80yIU1beH+DZoFMJ/3+3clMQb6CuGeVk
QESv0D+p7r4CVx3HYWcAbiFCveuxj8PfAaAtXvwAkgxyl6IHFp7lAPeUShnYnoh7hOK70PGqtOFL
fj30eTDgxtt69/uWn6+NPtKYhd5Y4j+OcAEJl1wltVvkOdd74g4PBcyKOw+uO9kx1EOH3CZI17wE
hSyS2ekFWVExjyvReyan0y7yaCbtmypbfG/znXVWkkcAW258ZdQKaYMS61q+oSq2hXibB6W615X2
3FxUlLWbakIHPLbiKoCm1MOgTzstX7F3Id6pzcIbrYB9x3LzIHc4+X+hHHG46SjNGOctaX49cTQ1
53XWrqovZoiUoOX0lhc8RL86vT4igVT/xM3xLc4B4s/N+DatxFVFY6tuLQ6GT3efqvK5wlA3cmFT
z8yJPDMNIFZD7RBuNr2goXZSHwPEaMEH71VuibKR4AvfROb4Xz0tIHVZJt3fQZTOa9Ql35c37NQA
BWuz9eMtRjU417i6fn5WmHYLSY1UrZyOWtZ+R3q7vWgPXOitfmZDfL6TvUxiZuvEe0ZbpF483wg9
OF6IMb+JKYlHG9ls0NJqmC06nQsIz6fmZC7NsOKqMv5M4S9sHfkbn1L/WryWDe1cN0BoQDspuGJ6
NFx+1m/aa1/z2Ff2pG9IARcJVuitli6tKndikjnu4LSVi8LeyTfxQ0hajMdJG0sfj7bhJU0dFx7q
u6z69mQSOBL7uXroV+6S59EP1bmPBasvM43C6OvSZOrNI+NLzpQytaV0bAIsQZ9Qp+Syy5I0C60n
6aU4MM3lvUbvRI6HLBVpvT78/qyzyhr6O0u219jiTGNJqvxvyrwfKBy5IDC53ljkfrZxlLpnnCxs
fCAT6R+9mRdQuBVqg0nVkCfsCdugnRylV2qU8i0iO9ywkTkf/mAfTdK6CwYI8X1Pxidr8hHbNcad
/8+mStTplnKMIKkWCSl+egeV4A/Ams31OsSdk4OdJ+FVZ6/Xl0HpV6nMtNbyhYrmKpimqFPelRVC
6Y7w2DMgZeUC5FNHIneeDlrQHGrprPWwabjHp+i8L12/1xngYVrEQRB6ARME49HWO4MIIMWeqfIi
mc7QG2tnlCkUDjgqPWA30sCLD9hjvfwxkT+S/NEjX2EoUHY9LxCZ3HxUfVKNbZgUYgawZryHk1Ur
tw4K+bIxWYbjE8El6jc4jh0u2AVJlRzj5h0vlj4qVd10mkhwUHgO6kIYffUM/fqZtrIEofsCY1lM
xS4SK1FOulZp+AilL1PgY1BeuzfkLIPkMaWTAF6YJ8njzvU5kkzZsvSQH1VHQwOcAdTOg9ou/Y5Q
NoQgko48aiAAAqyd70BIgw2HrN0Cx/0RLdyJNqv191j2Ias1AWX0d5adYVU2HpxSV3oXmtM1j2Lk
clmtbX6RnWCkcL5Xpa3tPVlLPmvWHv1Kca92vEmw/gNARU9Mc0YXM21XnGv2dMCbuOFbxiSN7/Mu
9/iON/WJUxMx1fXBbwS5oBvlRbz6Vb4Km/9zzzKBQwaolAj8XBQuy8hsbLNLoQjTZJWKemQ3Nw2O
X39yCJ2T4k7UZYHz977zOymnW/iE4Ja0fMUd5zrFH66+Qfl5Bp9N5lR4L8SqGEvyCXfNU1h0kA4c
Z9f8jUdYzRrAv5ZVTY0I6zkQkEIAmytrdDEokFCb2IDTb9vpXtYnbSWv1bUH5HdhAPVCcqH5tAwz
L4To5lZ8TL4dxbgCV6+gXULDBG5Pzwt0JoCse6/yiFz80Sz2VmLPT5mN2sXpWznytsQdNS7lG2fy
eRj3aS1BUqlG+dXAIVBtQU4BKk+1ApuykQaaFdPh28+bjHH95wc8vQSNEeKmTsb8XAGR7GZAP9Tq
wXRrpfiTOdN4+m9zgMnq7Zy0XixlRbn4hMDR9nCpZ3gFtaVqGzCdYIwHlpQqwPxUu/5uITuBuGgL
JPybrNTDse+l0xE0dPYb5Wutay7gzb7J4oMihdpsccli4zZcwDJBYPunCq6zyy5MaUkeRVIErUhp
dC5rWdKSC14xFP4gjm+OyEsvo1p4v5F3a6yHn37HFV0OuW0Hr+WFNt/JvCWIED+vBeUStfXIxLr5
wK7NPQC7KH7gDi2+RdtcLugnyjl6vnQdjCSgLT6kJ9vCGbniYODhTGdBZQYvnLZYmoUxuaPttVZk
52BRhWwZyQ99lhDcT9NuCR6/Gj2FuyjbkVdpdpymyc0XcEq5LI89pBoIl5tL2s6lKRjAnOgsT7mr
VmeUJ/EqXzbrJZ3V4sNFMMtltSm4hdkfMAMVyNA4GSmLJY7bqH9wiDPdZPj8/SoAVtwKps35ZxnA
Zsc5Pl9jqpvaKoLY9xBwWcsza5pPN+wr1WZp0MkwtgeVDBeB+Q17Vj4Eg9zR2cpWYVK3JGferDiV
fYjpLcnOJeM099iF1uFMZvNLTNnej7od+hgTpYpmMSsnYqc9t3IwG5ZgF+PLuh6HHN+LkWbsg9Te
7oPJYvht5ftBAVNre9uRJzE2LEDP85mv4/Ynlij5JjgSb1Fi7vf5aaQrp5X7eZ0JHsA0lC5hnGJt
N0oiEeWZc/hpl8q4OsqRPFnX64KCY/WnSOTQ3UgQCpbqoakJO1Ts7IFKFa4nXSIL3xAlocFKbYnp
2m0WN1H+uACO4/j3F/6qOUz8H3JcTFO68+kWse9cZd5c5dOD/OGR/7xxVHXiALZt9BEoOJCSi+lE
9nO50NRVcc7x+yiLzrfcn9wQUeWJK/G2mpNluMYjOVU8nfBRQzBPuhx6dDLnxMQZCRXsTYFgsoDS
PhE5WB82bToZOYQ3Oor8CCsR6rE/LJ95KWqberI/NW83drxguXfOMZ+aIT12vp5El2qSR/8PEO2I
Jh3A8cSjMoYZ6aHeK67xTLySdgFLHSYmciAztvDunY+pYcNiiupxhht0mvdJHHOCpq+y+Bxy72Dl
da5QXP0xYmDlbshr6suSfSZJnpYH7XLORN2M1yfwVegNJt5Izeiw7z5rdtwb/pVdmsRExQYRnKsR
IegghOOKSZafrIvVj2+0gVXhAShfF6J5f1uraeAX1pyRIqQ7iQsa9N4+Gy7O3f5AcEDoH336HEBt
xCddt9rTjyRpnHpsdYjDH5GFnG+9CCyRIi5Fyeq7xt7wHSKFRIRFErMBj9tKigdEnZtKrs7KAriT
p7eH146ZBbJXSHhFqVJJdef+XTgUYdhJodh4WAK1hGh9Hh/LD1+mnFpN062nXSG3Psz2Sn9MFqs2
DnPujZkd88tg789wviS3AbLp26vJoVUHkbL+uAoAtYhQWufO4wi7LAaOq+0sexDXjWs4ASYrJJ2c
VB2Ei11LE1wrKZ7JX5J4i0tTCuqP4cH4bx7dWiJrv83uG4Eud8JCH1N2NbQ0CyfZPQzcAq2Xwq7G
tdkM1QPpzzy7T/5zaFAry1DSaIbLWoBfwa+UPvp9/hpXDKTHENdH+KG08AhMj4TYPljcxWbDQfAz
ELtwzqZoAUi9aytRBNOQjFtaE/vNRPEsSaYK7FQ0vM7xVqink8oxxS0KeXxfMFtMKp8q0X7owXwV
1LsGXDvBEaw/J0gH4d5ydV9xhaoJ2lYd/9PqSS7J/yIaAiiwHomBif/DSKkP0gCe4mhqXgq/5+K9
qjDb//v9vfJFC6ciTOGsSjLT7xZYwCen3+mIOrnkmJqk0Ix9DLtvL6uQFtlk79uTjGvU1pqlTYVJ
j0iPr2Gbbz11KysTMVM1ruuIpziHTreFG4W7LPXod1ZAYzGwcZ+alu21siln3ksssWS+fcE3U1RY
4xJay95IbGQkOqwTD3Dbbrh6hRNUyrhupzW3qtEFlxDCYcAg+oXU2tuBJ77To/XcSXccfp9PjtwS
o/A7tRYcz6BJoO2xyy22F/3kyUsyOb5L1LSdmZlpsqw5Pa6OowdkcYeeUVqfGvj06SepLiRjOjmm
1VprZ+7NZaTzooY0NPfDfrTeW88YbVfofwNf+rIkJDmB7WHKj0pJmGamJje+LnpyKumWEFMV4r+Z
sVRRNuD9K5qplTzjn//BYCvNx/ZUUy3BPZ3+znjmccbqDdV6A896+4q9T967BHu9/KEkMcwhgMda
NtFrzGE2+8u7Ct60BatVYBr8YWb6BFx/fkXXZ8R4UHXvy6wJczzdYbqcr6m443EeXz/aJMZLWkgg
F1WtBdEkf9IzaYDnz2s5ZID9BOt77Ns9xsm/82Odp8nlOYCpnCeBvwW5xgZDifdGhNAiM9olumsp
Fdb/aMJf0BEfEq1Lk1G1uNJol/Zb+ZVlCiFrTHpunVPboQgFFM3fs3RiKJw4LUZuuzhYZoNqsshH
FkX9lRZqluW47dCIDtCY9l0BJdD26iaoa7rVDpScip58Rv9zhdZR4kItmn35fd+O1ysATcf/UMhK
aLFow5mhWLauFwbk86OqsijbyID6FTny0jQm5i994LoPMzy5PV/PuiXZT8Qu23ry1emdDXxVafYh
Xk7qq02QML3L2rmFDCAuTqBe/Sxk6QxNZsQw3BUOJlFMPA6N0FCNEOW9Si4thkuY1x06RGeBitZ+
mvYkLNkpWBvzf7PF3v8rqwd2RtsomVGshTWuidMslfaOfp2gaCRc5UoFu1+fZf+N2TU2UjCq0nXj
dUxdjR5G6tKPjxwB3OyplJgvJ5zj68iCM2gmTNa2bkH6oyLMzvg4wIljfbAUQiRSOvz1HTaL3Wjk
U/fuvpeoqFsHIdoKDATli50JUdZ+NMRQoiC5fTLy83DQ7xzYRxLx+2vHA5EKIDtWSXkkklsf4oII
CNsFz68Oe5fXC/Gslo4ChgKQDtjEcwWscXa63iB+1l7+FDsDhRNYkkyZ4IVBhzxEryeZc9xvmN0s
nCcvcahEiEg1oOpjSHRh7cAFbZ9kov5B4gpLTKpVLAVkfWGYyhf61L7soacE4Z+A4Bo8+n6WKFxm
ca0BXaoZFEgIh94Gv+5exKOUXYEBcFHwhYFjq2SO8nvVuPoZiFUsYeEw7p0VxtIsmmCidNj3uPCy
v89n9QBRSBPrGj4fQlJBqY3s+rnJ1uOk4ATYWUeQ0mWIuK4XWpoxvbVoo1+Tp/Ihlg8MIyKsiy+C
RX8WVPiexYdTOwhaWrlPTtA3bv+XO3nWy6zxGcZJ9o6Ejr8i/B7vi6Ca4/BKN3SFKPhVnPR3HEW/
BVGzCe1r/cSiUoH3U042VzbJmdTJVEDKjy4LAUmxXToyVLdOC5WpjSMX1DIgeSOSZvSgSZ4AeAzp
2zSsq5QI/cdo72WZJJbrk4XBPyU2nWLpYvQv/K2nXaX0Uw9ptpSoWeRcsfQHuvjvae7zw2q4eN/b
qJyZ2QuQFPnvQHHN3KN4VL7dEK+3gZpXqY/2amEf6VcG4IZxcxbRR6bH5+vSmi/Dp9c/W3uTZgYG
VagxbBr5XOJJkPxQUVqiIUjhQzxWc+okFAISQiyodsaXQ8XtFBB36Qv5lb2QJk9tmkBbPkhZ3EFq
26HZvigHZAXU7enes27nM+jDaKWM8FXusI/e6sLAtSi8svaSrjJFmk559tpf/+uYF0E6151Im6hA
mQERSApJVXG5/uTD4nKuCHGplpZ26ht7plKEBRrGhwY0hjwe2Dv7axScel7zQw8r2fUy1OXS0HhF
hh0ZbaLiQWAV7V5jNS+RSRBaOY00BzanxMhJSmKws76cqQw0T+a9oEid5lkw20q2bxn9JC2gt/t3
s8wihagAZ9rrSOG3ZmqGnxQATvQ54Pr2mU6PvMZa4MoTwItdymOeQpqTh73PdUNJBd2Yuqq6eDBj
6CSG7u8HBIu7c2xYN2e4ptdClMir/t7vl2iyPmXoDByEnsjfcCrl5JBFEDzNxWu6wKtgVvndsJBX
gCQuOWGECJ/cfQnEhZhK4sZfNkMKfvCiX/lasJbEZk4+AIxSfwzh30vgNqL4RlcZaZJKTVhe6RuM
JISilaPmMlIjSnLR7CpoupFAQU1UAMCYEsTL4KS3sXm/M+L3xazC6+pxIvZtcDuCC7Uv5bjyWq99
Y2lWBC1qX4y7ogfUgsZSQdJnU+6BotIv5aQSP/zKJjbr+MNHHUb3jFU4n7bkuNZM6GDhqlWM+ozq
HtPhfPrqFmjjoA974YmSpj51M6kk8jN5rFhWEhJn1wDZoWL0YJ72KLXev8o6ohSOWZUonPSdap7z
HYnwhKB/seyNup49GqqN+OEZyBqOab5H8Lhuo8P/cbHYt1olUqVc1ZZ3Nhb79XKowUo1YCKc3Q3D
VsTMtOswZDpa6u3BoYETEYjAy3JcE0K/9zDg1ZVuYUcjHNYau3r5vJNEv83hO0G4iaCfDXBDjJmp
xOTKYH2SInROLSOCK6yeSfcqQTqn5W0rgQ6hChiCdLHdjxM/pUkx5RutRjbzvUfrT2tkimw8O9mk
qM8Qw8i9KnbOpxLnn3Dq2r42DdZJM3jU/XB2lF1bPFMM+MxDr9Sr8AvxtycsvmLYfo+WfF5MK9qL
lrpSB8jCynIMCccgniZdgiZX6jgdOvUnr/UPIDku82V338Lr4p4XALVfXEvIBxvzpMgE9xNU2UQ8
+UocEA+0irg5SxDrvKcUSgeskB6/iOvRlK+Sn+nA7xvoXxPpS1H6QCkcYs4eBRyKMudEnLRwydnF
vYSXie59/CwIh2UkwzpOgTFjFhFkAbogecRS5gTnbOdAb8GnpymSaI/TGtNMJmIM2gQ8xD0pIVj0
Ta+kSqKX876SK4Q4MzflYguEy+wCu/xy8uP4LUArJadjBBd+rXT57kbPKPgCKgmc+zM+ItJTUHcA
JDN/dEv+se3aT6ze+Aid37ru0Y+tVt1OA+1hvu2Z0Tm8L1fMDEP7iHKFEj8K4xM1YJ+YKVgQQQwg
vnfZeI7InYtCWdsf55fJGRrhEzbKoZ711w+ikAZShQjqVUoethMdjavtiT+G9mUJlq/IwRHGhnj/
LfytWt36fYvAhlTdsmR9T5vp2Eh/Jcwpk2wSGrhXwVMV8u2WmgM00Bbx4i0jA83VymHubur/MjFb
JcHnkrgMRR03UOwLYgIJ1qPnmFVFDmrJ5istlBuAa8j20uHqeAyG12mwov5OK735uRczgGj8iSbw
oyMGcyc0MjoDIEKPy9xIyrxBYWhm+WtZk+78KIVQVTI8FCJe9pFR9bMC1TKr24ZqjLkKSFGmSHMm
3iu/4rCAP42sHJ/5n8mCoWT2QVLUCsVnbT2/D8I49jOvi4Zp1uxk2x/8xooCHfRO23n6CO1D1jGU
tXHkfdeM1DEUPcTASDaBPul4esnUfc8h3TYka/KOyVUZgx+I9AMNROk3NU1kOOIfUZerqFufHUZJ
rNE017k2YH2GtxKENMPpOUVFOFVeDwaZfN8PbDA68OTC94aPMPdsrKrzOViWlbbNmQ5XCy0DpBR6
IMDVJtFTs7MNiNN+j+U6ZWuGvg64cEb2hI0ko2g7p2xrA93BjsypFbEFqLtaFV2pdChmq4FBwMbi
ikziJa0hFZ5SYMNLv3hGt4VOQLfylZKkVNz4W1AzSc50AQ55tQTHr5kBiAyF14FcIMONAvClevnA
OTpEb+0j/toPsgbHxgrhseVqT2EqzCiWJDiWIRn5JBRnLvzDV0C05YnLNhmr3Ap8vL8sxl7j2tpH
9C7ReUtJz543N19sgXQOLeWYwgRePEwV8iWMrl3v5RcONsumiH7GNAPv2hWrXFN6EVPIFnlZgHTc
Ok8rNbOF0CsQtA6ujmQ9HovLwEWAaU685f3hilb4l7/byGT2JAieCp3bji9jpG4xzecVKaiNbZy/
wwBCDnKKXwy6gT/cibkOQZTCYu+CxbOi9YSd1v45Qa4BWu7IOXeOONzvx3njRrQabiam+qfxB8Ac
VhSzjLMSm3ER7pHip01GiV1rcK3s/4KvJUrbEvifuzaXRK+dmT4KRMHPbkfJmmt1Ie3Tx46eRVND
lO7l+Iij6dZg/Akqt/VgEKL9s1YahUJH8nV2z1G6TD8O6Rdtmhdxby9FSlpl8CqQKOvP5/9nxzK3
e/nahA/k06w7TpPk/MwJO4eYw8QVzFjsPaHmrCRRY22ybx7dcz6eY07lYioF+zDjpa6uaaMiGiDB
bwXJerHa6A/6Rd217A8jdWtEGeioZjfxQ/jV5U4Y/o2tneeoXEaz9wm/NCqqfT2wSrnROabpRfGf
TjIrT3WmjhmM0+zXXmSfiJczJUlOcwxHqzQK69GCpuQcQLuLA/IqZXUJPSkWq4Hc5FgvFaH3c+hR
fIxw1Xo1fhgrZVSsj+3sTW767JiU7YF/h8AJ2PBncmAr1L45yUkCvSSq9+u1uOt4giw3nLLj/u0F
R1XW8DVrMF3x7wx9p1vw3GX2P2HDQoE3uxA3+a0+EsDnRcdMtobyxlX60NzN+rZCL1ckHcJUQCjU
VHXRapkzbRhv6sqxDScQWEz+MC0haToIInFBg8z2M+3L5EYBzLBc9i8df0RJqENPPWVOBeNIPcXk
oDFWuqHsZXT+OM/Q++hWiGvGRHY07AMdty7PlU/xOgbaxPwut1BI+MmCCiW6BRElMVSVWOX/uFhl
DKRZm5ZzN4VJXkx+/Ijd2CpWtq7r5mxa7rR3vbXxPa5Q3/Tod8AL3C357kT+Lsao+ISqqC7SSg/J
iKd2BFtN/5l6WVJy8i3ptzNlE1ywoYvQ2TWjaOSzBppSRTNV9o2j2g0/1ocxt3luVOFKS9f9f3fZ
lXOLAvulpUW1ImYW7kKtBdsVidZDNuQFsCX1YCXzYil2bvEXpO8Wwagc/0fjXYd1nyopSnyPSHg2
4D2Cq418NZ/Rzo+ordAF2cqWRLsPyTTlFfZCWTTdi4GEi+OcwB0gqUjdGlFauzgXmZ0TnDeqDTY9
triDVfc/zJPsUAw8ckqmIeMGmCOZlSsnXgh7AOfJM8MBnzQf+6+J17ZwanMO43fVRAfO+h/lq3Mm
OfAsK1/70t4iPJcrUtLELzwB7KODm9H+fdG//R/iT9HxcCT5Ed1H2huqpyckAJcRL2wjgHuXnkFJ
C+swf+f/H87xMk8Ahw16LvCus1M77Puqc9aUN9UJWfc5b2PGNdJocMZ/DxaTZSklV6gCiQfJRFpP
9BBwabFWRP3JicDoydubrQm3bZz/fgrDq6TMhvMVXoeDt+029Se4ApKQfZPhyVJMwnyaWUFGkof8
UdfQWkjNpom1VsMN9/sI+TpHX0cCogPvrnTMDNc+Y/nP62+7wyJo/tOuDYUAvC6EHzHhYtQmugIv
4xkf/u2DT4opuFItlxpCW81W1oPrGaq65575CM/xEXEaU6+WM8AeKPxwS1Vw+iBYptKtkvI/sqDO
9Z4q7RR1Uu6GuMwr+9MOa8fWwKBp2IeNDTG0texH5r9s3B5AF3NS4QKX/7LbGiciEQXZGQuCKLaa
w3HlPI6wfcKVHI8dK3OUN3h2rP5OR3xacjNdaClibGjcei+G2WNbvDeNSJlu7cTtZwAkC+y6aLm1
e8AcFrcLBUP3fxZNI7cf9mTVMU3/g5a7cXGl+duYaPaIH5GyAEDR8xrPKbJmnFXa+vjujARFnv9F
o/D9dQp0R5i/3bk4oAdIfQGy5031fxT9djM4Q0rqdRe8IEEvGfl0aDBPRFwAznqRi+PYeVyYhdIx
jQgVcnn2Ov04ZC3SPHCHOiWwdvSb1zwMe25vgko9el9WCs4drs5xDPxTaXt2MQQh/EX8ySRtyz8T
u72L1BxwmduV1zA2veuNR8an2RCPuVE9BVTHDFQH9zEiuC6qI2fwCNrRH9pZ97Ym0jlDzi6tKUWm
izcv5VwkfBxtor+tKC2c4tzCgS6xHSsX8BE8+U4r2Ny3Q49rySqrW4AUJkcmMKrin/AWaBVyXf3D
zuGvjQE8hreXCaHvvqMPMJ8U2LXj4pBWUX7xq418d7Ey3tg5IlUUo8LcZXHQc1NZKqmtt4OsQupW
4jLx3mFNkkFnmvB5Me73IZt0tQusZ6hZ5cTjfFe7KkLlXet3WLUXEUoGuNuXkelKNSrUJZoEWjam
gPhxDiF6Q05pr1i0TNd8IZ2PwK+6ff7ZBRACTx5/WDzdrCGNsvgH8699gmR1NDPxxrV60hpDSi0S
bfPeUJWHy63zTgXoxH4ayGREuhTCKsnT3EjMde7U7SNF1gtfehBEJDsut9du6l5vIw3951AUI0bi
jLQWOnFEJxjMdpwCryir4Ep7GkYcbdHFX1hFx7J5nIhfz4ANwC6HoUVeWHbpYK2/9YTNHGNxJ3KZ
nycbbaAdTpbkcPnXMU6ZMqm4X93r+sNc3Ui7QG2+c8dz+e73ljq9pjEzSfpEkFXzEEatSyzfOfxo
VNDPBy/Bh6QVRIvZfIo897Wqp5phn6/8vumx1zMPTcbTIATD0hMS7l+GcaERdGZrpAv2Ak7t4j6Z
8VA/yxAXLfRbNc9mUXlyEpt/Jp1IqbhdTdDM4uUxp5adbENEVHwMsixn3gD3WfvfrJi/2KUs9EMH
G92OCDKb66KYzI3gQegp/7aMtZzV2ovSXjtvSoDaLemENFZ/MyHfzGYGhkxgOS0sUc/xXwPBgSjS
bUgh58cWkGGst06ansNQ5ipsG/Kg9VIPR8iU2mFXH7XXeoRUlHv677gn1mxxqnXwo13BtkpeaC9d
dQxaj4NLf9BglBlti1dMuOpV4O6Cp+sXaddRMvOxocG9S/h+5wilXCVt4AuaBeBa/Gm7BYWw2Qx4
uvZ8nVRkGW5UVa0eIrc2ebwuvCn+0WOvBr1k8VXg4yhgVyD2gnECRSXkmtfDxRqrxFaGtgnFXStU
eEDQAx/XQDx4llDASE7uMg9zQjfZz5J0kTo8NLlo5rDuT7+PmP5uXfxJ0ovUhgXghsDYC0dXRQdl
uvcvdX/EUJf2qWydoZ/uS/NnM8mOTty9kSRZQELStx+nHgGhnY097AfjKH0m/KdMbqfUKR5CITHB
n6nyAfcqUppk4sAOos2WnXaeK7P33QHHsOvdIkM1okfUrXy98FnuvwsnhqZbITAWGo2I4CHDunKL
OPuz6T8UW2Ier1RjsQ8hS7iaZniRhRQX3/OHI99Q1D+dDW/VQdd93pkZXt8JvYY4lE2RZeZHvLTY
LbVjdwMoidLzFfzCKLk7Un4GVlPQOeqtU0VKmbtE5Alk/yCTRtsi9OPbh2dPRY6Zcr8nS3JgIMPU
S9O8+ICo4PkTVkPtd/cXijKqt0Le6gILrcbl9faMjh0cbuM9Zy3DyMsP9tuW2nlp/tBQMVqtkx/Z
wF/1rUHhLvJmTA8zmltUPLAre5pMfPEQskvmYAqZ5w4PcXwNl8iB2FQnIwqyGh5P0+QJNqo8Up8w
wO0H45/alrZYCC7B+Oe9huK7vSIKCmpYzUI/McvGXlweV1Pl6l5bdJbYbhBVZlHRys/Y61VuCzDH
yB9lV5T/+GKljABJvc0ZL6o8xovZNFmUWMu3/b1N9h0sZNbFLlUoAdTaET60A4cd65D717DYMBKo
mqKLBtt26RgDZ3gne3Wvs5zZ+UEy/T5FXmcH7+dYavOZRyG3Pya2tRXfZtzrxhN6nL3fk3JQ/ygE
bgBJYiH4vqo7tiHqVbMNmDs/cwVAQ8QM/DMAtfeqxDrHjF4jREzfWzGBLCc2Q+mdkmH8pv4ruTip
P10hc7lSzXaWcrLD2NNOtMPGyPKN420UotXrA+a2P4haUW0/zB4TsUBWFdX5Uyl77zHlePX+pFBA
HefbMLzf07Nej0hwoJDUrTCAqeGDJkV6QmipuRsFYJAGFfkGTqqSgCwOxZqhgi8O8VO3vIX4Ntrk
o2ezrkMl/MxecDUlzVKEE7zDhyM5BMd5zlWkhbMnroG10PhF8o5A8+ci6y9YTAdKfgEWY/q5mDk/
Jupv3sgjXVzclC+vmFncwztervGkPhnOWlpe3SoxAMJOtBR92YeKFUWN/p+FSJTDlIt82xg7qsp4
iXrJHcBuVpsE6yhFEkilTNw/7fNQqIu2J+ww9pRAVSwJvj+jzuHm1kRx2l2aLdYHg/H3z6aHc4om
wVPj6sz2vyZkYUfCWLzWF68iI8BGS7/B/zmrHaoVKmVvJlHofFl487RP1sa9VVi2RSAyXcqvtUzE
f2SzMHZ3GLqrT6Adw04N9/gvycjXJSAPtSPxD0BeK2seTYFiLv6JPSmTLjS3yAZ8aiTrzZ2z9L1S
sbqRQ8Vxmp/98mBZvvgNPPd0ZwhvJtIQ5UVBkkznROerRMiaYuos7cOx50caJFKIBvi5WtiBx330
RU0//l7xxF4RE6nbbQ/ACWsTBaF/fUdDVUZTFnETx9Cs/1E0bmiiDRYWrkYltYTdUemv+hca0Dys
/vi/dKA0lNrJUVITsNC+LibLC+YayizVVNswQi3eBQq7fKUACqG9UBc1azVgg5FwEEfMTtRr5jAP
aZs90a0puxIvRh6cB59T9NFlBJrw4JugHleYIJan5SercnXz89wZDfWDXQQtXouOoIkP/VmgzOOW
LA1BwLyZXHp/A6mFQuuaAdXDwGTGLUgEWVRGyn2Aj/y9kABx6HDCbqjBJZ2LDfeNqQwOYWYPEfpO
V4amYoJvIDp0kzUGByrK+PtX5H3taOxYbMxWPYKCY2qNQUfT9ze4odiZKUUqqERpNVioiSwj7JEH
DVFLHEC154TB9BLDnK0smPBZqpg8Sdeu9QDC3XzPSfJhPrNx/InXsQ0gAmsEY/bCIU69NzxMdWPd
vyAGcwNywfArxcT5XGukVM7INboYLZByXOR2EfakURUZac4PXRalOMyuffeHA7T8Ke1syGalCUQ5
Qsf8LKRzRJEAasP8QBuYcaUiuNpJV+8imZs+rR40PkfVfuE26047Q5BVTF0NX6xevR3WtuH1IJ2i
ybwQZE8qNDTE5kH6T+M4qpwA6eaXCGnir5q2J1YWrlJxVt/uaWM1QEbt+kP9ODfCmgpQ+j3Z1Iyp
MdZpwxRx9aA5lKDSV8O269OMF5WSaskrWoD2tDFMExUyPuZrdThgYsjhz2LNhzYZtB52kxp05UmQ
mskBVu0zwSqQXF8y3xK3c1Mya8mFB+tKZfbUjGI2z7lo8i3dEuORtDPUqPjiSkShltSVPW6X2232
A4camAi2RVzpZMZUqhNpUcR7Ml0fBsPh/LML1TvUn7eAxq6J3P0hRHNtLqujpLc178UX2Trmgnge
vrY1xVHlI7ZkWvu9lBJZrh+CASTIUFrv5inLquAP+d8IPn/CvwIdjCYYje3Bj5xfVzBepruSLf2C
dLoguxsh37j0ZLtDQl1Y19JtjyqkUIBs7DkgTWB+XVe8ILJXZR99LKWQC1gHbS1BnrE37nmBpOHp
vgv9fowpsaNgIyhJ3uWZBruTDwbJtzsOpC+7kVycqleTTzIvGCUx522/qn5d7HkOiTYWzgFy4j/N
FHPcM50puCSMT23bJy/bRLYrsb9+C2r1lwQf2/Q29UFeX6+OlYrPfP/bMWejJkgSjCsXBsV1/c2a
L+qmnsPF5EaOL9UeQgA0ouK1/FZqwuymy3QJR8LNdYjiLgKkh/afl87r7hemovVyEhfbZtt0ynKP
pasTCU0j/Sm7h23MEZO/dHEr5cKM+89FvPeyxO8FqaGI5xj5BtYsCxTyEsynw5Xh+JWyiRf0Gdz3
SDClXTbE6szvj2Ea5AEacjpCNdSA/xlahrKnapWEr4CGm/Qu4DyQNtN60zPwhIVrzfEmBPs87UHE
p1EALpLMcpOQ++LAdGSQMHpfmxzrCVOgUyEg1PHTX/9ELEvAYZfty49svhsOya7GO/eGmomm6c4v
HTX/weefViKRnpt69XNEso0ZNbTxgAoupTUZ+qQB6xdQNaJuakTn/Js54xYg23ngaxHw44EK9lJz
R+wOpXsaDdnI/Endkv+8/js7inp312gUAH8gEzuhpKp7DBSonpPF8XtVqdam4Ddwk2H0MNiFyHHq
FEnuusjapl44xnJaNqZGsswMRTsT+4XsLR/kDbfKHgdp+QZ8kfjJmOeO0vyMVHIlBuMsLBMe9rLZ
YIHZ2XI93i8o7m5St+z/KmXVmKlNJMM5Gx5HVH63+SoISqcfe2pUXrTXikrLuDVnfKlfIDdGRg74
h9AAvA7Hp3rUSoeYdsJCD8YiZGn2RU75Jea4E9qOcNMXo+h0Ls82R8y/VKI/lWKG5mYPzabaNNgx
D2EsqIJzImtS2MPHWAgHDcL9kjIP6592dftqpSDlHnJXSeNToVTehAoZxTpt6LNUDRAGac+RkeEr
bRArzm+1/ldS1y2CDwBtkfB84Me5zYBqaeEb5vtvqwRNtKNjeTxX1+LeZlisgXX3lfXBXCOI6jXs
Y1UmZXlcN4M2utSg9ZmkXekukqBRu+W7+SZmG6haYxVd5EzwdrUKg029eNmcljJTV6xgn39CMrhd
2IYpdbqbkVk6kg07kz6m2xGngRF7Url38seDuA9m+CVsHac647T/6QL5yA0Ah/6MopHjvxsVhZLe
j9nkiXdx9V5aMpPxzR3Xbjm6tUFpEtofMMsj7t3yPG89El+8uL1+nU0AtWbl9tfr09TgbXVG+4al
NAKt3Rp3XJie7OE9i3VBtOAUceiSMO8MuS/8KLSKvmx3OEv3NTkuTYX3QBQHQJFiwlDXtviIXCNV
GviojglvjHqrHLLTTu3wQa5Bfwg9NgJm4ZS+JRE3L2Lx93vxOhnq13xAqPNW3sOPvnjSD77skaL1
2PHkxWgViOoLtHQ3ETa6nXBjrGB18O1TgJgIHtDXXJaLWyFrp0BlzyxnZHPqTIOGAErBIJsvDIsv
DXWr+8oDjfu7A+0wE4/n07juT9RUt4HacbxA1Pt/Sw7y6/apaEJTOpNKcOIsommDuN7bjZME8vlD
tzKdZ9+3DIg3LbvJNIK7I/kf8ONqzoTeIijtY4TqWsGKXai3kzrDteOtiRzh78N+pcRtfsZz9vET
JxJjN6QwGkQCbsPPBGRWyS74iLM9unRK7vb5WAMbZTOHyyf2YE9VBSM68Bzv8+JgYV54FR3YMbCF
EtYtdM1al8EtcX+KP1Y0+xC+dazUXivjXC62NS9Ut8C4/1E/r20BAYoKCY3GTLERBFwEEUQ96AKq
4ykcfCtywl58T5e1Xc9r6IYR78c/IvIUcmaiAtxt9t0S/0V5IAjNZ76CIGMrDPxa7lgwGTuoqG6Q
jyTnAlYlQSXmNdhGVZGefn/wNOTLG2H/KXw4VWKxkPPlHyzP78afspLBmfwggCz+yWlq1vxnF4Yq
+P8A7ynCOtCv7EyMVCLcQ7SmbqPkbdq+UARltdueUoNCGkJXJoIKAgf37NY1jhJfGoCLo/Gd5Y/y
hPgMbLB7hun4flg7aCX2wZ2TmWDcuNOzaJ+m3kotru/lA1naKlfSgJxvk8rvBEt29CTbbtJ8LCj4
TfTlmDxIzUkcOsaGqfCB8V3hFStqsBqzvsGp8+0QyElD8QYe4mnKf4hOzUEyffTdBBjaLg5Qm49L
z6OoC2n74gUPYEKpPc8MGod4Yyc3pn8dNBktaxe7KbesuOVpJiVsRpoYQLXzsCbIqbjv7xRmKzFQ
dwnUktGDFwkA09IG/gPveVV9jOCtyDF7UztgACd1+0crfUwhbHS6DDYtenSZMdvy9WTe8bgSFMDG
CISizK1EUFtlDe5IMjZOTOU6ml6whsE9QvursuHaXuVFmMMCPZreVE0d0bfHq7V3cXiHw2/nNNaj
kh3cduxPpvndVHjHtMA/4EtUQWKAYgqOjSM+PdowMT4/sdcOWNfpbNR0qyw+tlmJe22Z+XvhiMP3
eNa3sC/KYUADmMuVVxX35ZlHITBejrMrgpnyhv8CG+KWVqvvC7DBEA0tn9mAkMF5bpPVbZZEYT4H
cYEqVUZIONPc8FSIURuOWDUyIT3I6PbUwXRudrwpshX1AazuRX9prQWxVYGs+hkUZVI9leZmBoig
0RT1BLqw5Ol6EoKj6mv/k7yGMaLOnpvlacfRL31LDkmfb9uOIpGJ6Nhi17p/01aUHNEnqvYPGZLX
CjWhUDNKGYBq0a20LyzPkdiE5UDcXBLK33WieGTLaGvSUI6vlG+eGUJ8HyhckuuPXas2IzTlivSt
Q0IVJxb0J20Lo+nXGERfD+vc5HNWq5vw2zNCYyDxKT4f5qSCewXAT7z3/xc7F9ZPz9b+N9RK4zQi
Oc0ZgNZ5XEG/HSe8cwhkm9gU9uPJW7LZourACBEpNmqdxv40wq37ODzH6FCR32CeKN021U83MMw3
BJzdbz0h9AAcf9RYhL66rsiFIaJ0eCc5LLwAFsGJhiKYrVUwAJ/2DOsi4fjbYHlN//rQy5ZyuYY9
doC7GLYPzd3KiF69XJ4JLfBAehnjXZlXKi25x0ielWO9/AQmG2Ws5mU9+KoO81xGnQ5rmYcOYaEn
hQ3GfDvT20wwmlp1WkTWFNnasYx4bSIa1o3HMF1CZAJgBn9VKgCSmMdcN/kd4me8KxyWPJEpubdm
aKfPCtYTFvMyL7Rp/Yy5dmSG0aKuyYsxGA1MwCzyylZPlnenbcu9E9CYB86eb6+sBIxht1BTWyDP
bKp2OHG/pz8DHCMq824zDr58Qd9XEwJFiP1Q7BudMpaQnMLDjb6jz9I54VGzEGWeXffGjw7jjnIq
u3ZyJZHVetgj8TZYlOShiE+a3nMzxIm0cl8sj+JLdawkJdQkJj9b5O63ucl13toYmPGRg/Lfufjb
sMxqHWibWOIoWfhB/BOAwzH3sdJZKAqM239aL8MgdZ6GZerJfQbPjTGN9AftIRX9mq8jpSe9qXao
IPmcTOn4R/2NhIw2kRUObna6A0pyMwnu/ZfMZume5/B26kTEYjYJ/MEswBxtUz+o8Q/l6SxeLtku
5ZKQ9EropPcFqjKwMIVYFu50s4M9guPM6/hIpDer+5LSLocQCFDwYWN+TeAcOTu1SXI0iw8hN9b2
hT02aSuqZiNgsNUqaYadTSjnFfLeWEb7fUpWgNr9iOmEn/xydtH7MlH5oK8KzDUWTo8xQoerQ6UL
FlRF7WNUb22b0xyzT9NUMxkjdzrTLF6fxC4YuDikDVYHaugnrJVP2Cw3BJVWMmN43gN5hzmmhPdv
kgSGZGVOprVntO5wY4cRX8K0vfC3uQkjwqM10R+aEIpktCJSysrOG2HAnAVA8O0oG733LbyCfs6Q
r0VJTd4lVRjlEZcx/cVN0ai9fZrUNcwCfHxfHsoENfO27moutoN65XnaAneBbvh6jfsr0hexw0SO
yAOWkFAYk/MzNeqzab7Krq1Ix5NF8ioEbPGMjwlLfC11poOPBkgmAdcTO6I0rV9sTD2QYkjDnsgJ
09H6vHLgy+45LPe31Mn8ueSqLfxUHlRySc0Q9IAWWvweZDkjDE7/yVNXRQ1XMvQTJPA8MAurjU0M
hmw3GtAiel7VF6WexTRzX8Hw2XSRKvOgYyt7C7pUVvUUTupq5NpRS2BBgO/dzfwrFjOzQ6a5c6MV
pseARhLgrhzh3uvAKFnjbFLIIsY5v+b76RGCAp/j3waYevxBY78lzukrvUGWX+AuHG0NWYISR+BU
zJ9UnO60A4ZUcR9S+oN9VOx1l99lEgZWbkYdAZhWCOgICPgQkVVBnRb5oD8b08/6dB4ffMy7xYro
zi8tJQJCpq2WVDTnxdMq8/H2mfqLTJNDTwflfL9ku2pSl0UoCeKO72dJaCRydUaCaQjnaetX7s+T
cfyj3/C9Q8mEORVNsoTb4oIdDkcFNsOFkL0fJ9FH6M5lDG/gDOAOgWaTFa+XfKVYXloKWqDXK+mt
0T8CuIJn+xCk4WPjIIHblRD4X/UzCgDQGI+IUlw/pXSI3ImvVwI9vwB8s7MhDvcl1hBj5McdfiEN
l8B7bIlSGFOGLXa6iHMj4qGJWDzbgPAq75206OepCMmCoX1WB5ZFjKLyI/2ayxe0QztQh9Q05wCz
csPHIpuK+uumkw+K9gluFALVUQlXVvQwtHQV95qPSqu8oL+BUT+gv0foJi8C+U4NkF5SezrKtFNy
XBNIfAeP0FaGgNZhMG7Onz8sD5AXwJiKEVrnRn1WzN8bdcogR/YV4l/QUIX98C9WyV+bAdArtj0C
IQFBzuPxcfO+JBLwuW2sIxBYbq1wD5A5gZaDXK5hy6jdEK5rl6+5uJy97RIJVnRVSxeYOzsoSj5O
60Z2j6mxgqOyksUN0ervKaknIU0HDYp5dxfcDffRKpSH8JyBQczg149ekuVepbKht06vmRB1WaNU
OAtLpuij7tkemDA7T1O0YCqRxL65UbhZ282m30yY4dLGjbOIe8lJvTjNMId3gBPistOrLgTOZu3U
v+x+wLEP0DWnDy7P1IDy18sZBbbFJMbUydXOHOwTcehFgqCjufHZ+AgHQo48exyn1/GfzkACGwD+
VpoNdPuQmxSmI1uo9Dd9sPKzt6Rk45vY+rj1Tmg6TJYHGCx5QKuUVASIVS5uAZFVJVPvBq9LZS3w
1p7eZoFIJj6JkWOPHMZnRoLJICc37rB+BywfMvj9dGASLP2ij/CjpOtMY2oGgmY/dkJMY+EubJYx
hmtDjcZW31cU3wF2Kq/Vt+X7GVBdz4r/ZICROQMMzba77V2/BgEOmL1Nwd0BNYJHxohlFP9tgt9C
Ze88HfWTKSjNlAbniNfZ0dWhS1uUpYC3i0NgCJ3AXyH7Auw8rkFi2ZfQUdGiqWIanZMR34vvc8en
bMPaFx1J44hKw+n3fNYbomc8MXQFYBze8BkQuZckN88Jjm7NjmcS0FM6FRVlEIjdwV9jwP+y9iuT
JN944rKbzrp0zHoXueTpFDsAvnZQi6CucxeocPUP6A4FL/5BE4d3qAQF9XSMlxZzOwJvRjX8IeSP
lGGm4WoXAPeccrK9qJ1HgTjThhL0XrvJTKt2Lpv5muFarbD5y6rsUCxS17XJNECPFEVnPI71hk7s
aN5jldEKXMbxo3qEjifZlfcZwmpjqNHghVRmBm8gLt5KGc71ORd01zaVv/4zRnZwg3xIShsiZFeO
Dhoy5Zw8WXZFUSGbXeyG4RAPUeAPTeo3rQvvo1zvC0D3yIOzRrvEDSvddGjV4hzbdofIQUvO7bDg
sR8+KD8cgkm5Q6+P4K2GcbMJ+Pb8QOs33PAZm0xPC/GQuSZGspBAvMplFWU6P/YZ2eA/drKfV5dP
Sqosd8H1TigraCUw5pSdfdojYbpN7Vn3i8Vb5M8hNW+8j9hofUDHgQrPtOziMT+Bvo7UDEA8N6WN
hL/uhJpkeRzGnJXYd+mp8isU+XWhGKyLZJ7jRDUapeITSFeOIaXZLRvTkPIDvsteOmZVmVDTBBPb
aFTYQ045DsWzZ/jCT5bEgxLYHq/r0Sz+w3F7OWI0fvDFYugUSLCZKccWHUx6vWbt+a3Wy+xbr2Fp
T+uWFDjUX4oChOXkLJdxsYpxwt2vJGhGhAuh5ZOxb4xCHFvtgrdv4ShMxhI16dcdS0ZOpmsR+yWz
Giwp4bEpQUhZKoSyYNrCRjKVK11LdhsaYOec3HpHZp5SCefjGSE9F1gumfMJrIQ+xPFi6xojrmuj
sN19c+QOYjf3IIXCrKzzRS5HBWXIlMYY+FTuyba4zNxVmFMNyQoAUKWAU0Qed0Lh2D3MQjwNbeJn
2z4lwLNEF6aQvsDwk/aBYQ3pFxeKS+ELXZRjqjwlGSAI1kWKg72XAtObogADMiCJ7vWkYbDGq5Sn
VSrvK0pVzOq+UphTJEK8I5J/qo+SvIuFUaaRhSxt3GNTuf2IRKuVE5hzCjLOtiAWHy25KjuslNaW
05DCr+30aG4iaOYgcGNeYhox24mPnfMS9DOejCbv5DlSG5q8KioU15ulhu6nxzn59Fulv0x4Te5F
CltIfbBQHzwbfADaW4dEx1/WrckJhkBQoSTrPO0OMgdxJK4E57xe+Z2v8I3p3oYHksjyhSPPHxxB
jDUKUxzgUX8lZK09EtfZZtjAOnV5XHrkX4PPcixAmcgy23IBAsJm7Haqnw1wqUhFDuQHCsd4MA5O
V83J4GhsbaXHl2fEJlYL5zevmpgX7gU7bCdMJrznuIm4clkqUMWaXJSPhcyvNMkiJyeKuNRXukO/
a9/FKmN6F85Qx4kote7l0jioa8p1x/TP+j2lilyKZ/xm0qSbgZDmqTMH51PjhUIFGgiSGKUAipVB
tCxyNpQqT1SNaMIYj9fZpjh6EAlDAM12yj4fzrLUeppChu+dMTz9RfKdqA95QdwlXjOF3vfNQJ8u
MyYepwDNoJl0oJEI9Qqdo0UN7Rc4SXlolp9UyLoDzbDH78L5UqIbgu/Zowh7zpXIljovUmSPKuEw
FwId3ns+D5Z1XunOtHjWmxKbhjGoO0XQ9SIkm+uLQU0Vv03sAtZJMML/D5Fpfgl1m0gloLUWs44V
3ly0PiLxPS2PcixPJQuPAcAZh8pJ9ArHBW9HZkepWBNbfoX8SVOmBc09KmoJ350zpfXIWn4OL3hN
k39XxO1SMGk3bFmNalKKqn/ddZ3Hk5/QvWXZqIv4rmtnhH6zQpvaYEGBeCjuePK5mHF1Ncdma+h5
8UiA2jWIYZyOrWrE1n8UtZW6ViZogEhnRjbSobWZNRf5Ue7UWXVFYQjnqbhhmupzmyZ+xJY20qf2
xVK85ggDcJEvW5HnGWfp9p8vVpIsZRv7by1/ka/jqlX5virWSApnFEjNo2Cl9op1fWWtBoZvVexX
Bnn+WDZf+NW4Yo4BRJchdqC8oSAKNVU1ooYfY4nHD4nJG/dd08kZq70OGGjs9Un59AVECq93vdBr
218ptuE91rTZHxt1ETVdlkysKJjcOgrlFx6s6I9DzAgoReP743T3Kl+nFtKzwb/v7EOdreac6+u7
C2WYWFNwzTMeVd/aszI3zJx0u9zn9ekQmwyj/+WCIEMeVtWRBYWy11Tsvo8tkkN+lUQeSWcluZ0B
g+KEpMKO9CFCwSICuZPLPoHnPVRMLdyGTnCFIs3DKejJaS/9EN1DY3ulfcxibleHQBHVqhxCaJk2
STw17KypIhciRemJykVkRt6kU/JxpEqZg5QU6xzYJN3ICqyp74m8v3qux2XXew85SGuexxHwj47R
oHlmZsp8OF+lZqtsIJraky1rQhl9QA/uDTAbNnj0Hz+rNrtmynykFocmU3uFBSGxwZZ3QlYEht4D
lA4cusjwsQmCwnmyoaQvsGHWd6xq1VbuoKd6cpa9oSG/+PlMqn7vs9F0kSYqYy/6BkLs9NoVo8/2
9AaQdTieV2iC6mhW80KZX8Ib+ipAtRhi8ZvNksqAwUJjWCleUvYaIDHrnC8KnaAxkI4LtcC7w0Sa
eL0VcpgTiHS8O8cg44sgajhodD+6ePa83IM3jpdb/miZLz9UQlRq1WZdQYGgq5DHkyGocE5/seDQ
e53T5kQG8P3qr3x8r9c5bL+R+Yrnvm1G5Iv3fO7lyQrWCQtPsZIsIab4xcbp3X0SlJJVriBoVEnh
1aCmlbp64DrsCkC0P4f3z+ifdo+qk3CvhPwJwkdMrsQAq7jGVTGA3Rz7vnHuAmRZXlhD9effV3gB
JScYNvdSKuGkA5y72Se/64HzImYsdokEEdqaUcC/8BbjDV55aSkQQF10qzpjF784k5SwEkInOZQJ
xF8B6vLcIKphQK3/7wBKXynUdZsT08YIg7Ieh3i6AkKOg4XEikPwzkVFW5CFQfpirlCaGuZKX1aH
XmAFtUom3dtxwzkIe4kiBD7aMxCq1ECf+twoi0aK0Pv0aFMCzkf5mdAJu5RcjCFt4jyvGvfFmwd4
AIUYjmBQDUDyUSFvIvVidlsZa8QAA+8F5bDEl9C4QUwFn3pdfMtWTu8V+gMCgk+TbQiV/p3F+1sd
c3s49CUC19Z+NjxF6g7vWc0C5EXmFZ+saq286aipkRu/9FSQdNNKW5NEjvJRkxsBlSfV8e2aTLGS
Bx3Z5DlKpurBhwPOISNEhKmJf+JNwUStgdFOqNUAi0lr+6OKBKR/jvtaxqDYwJEnDogNv+3bFvve
pHWRIMGJtVHMUPshCCNG0C1CwVy3haAgW/O6gi1Cn253srgXF58FzSrJQugelETgztqrPK+l8VgG
AZ5V+ujxUSx3dFmpxMv+7DN40aydVsoCSxM04yYurV6Lc/As0EyoRlpnYMeQgrCZfTrh7abSq3pL
jtWd7Pqqdzyq2Q+kbilSgVfbkDMhfM3e0pQkmna0W9dUCIdJjIKIjivqZ0M2DKB5ygdH6yBmOQ/s
vdwPVuvN/AWCIOiZvq2KUmukeuf+kDkw3NL9ATyX6wXFKvikbmbjY6S1modhAuszdwWNWLLDTOHo
YM4tYqXD/aBo/iJ3rrTaCv6y7KOTv9ua5oCnat8GTZ3y8rXExufLCNzgFBw4PAUXBb9gNziWEXpS
v3qOi8T6Ghc1gg26HTuBFIEGGq02R6LUVYXvfgcnpmAJK/i/XO/pXIBIbCqiE6WvGUn1Mlq6DBsM
SobJAXdKE0AnU58kxIdELq5O/Ri38EpHaElGGnxa02Q8YVXwQIg8kURvZdJyuvX/9dlAeefmpZF5
ac8JR/Hckt9Ipp6qo8GX2R3dtB2FcEXzUIlJWxujwdKrwTM1YtGns2z0P7X3GZIr1CwIIxBAUqlR
eADIJVgFKkP0JbQ/9UOlEzAtpTnGmStnl1IzJ7UJwsJv+Mm5IRGF7wRDO3k4RK97B0XzahLlrvLv
KTHaF8s3IFcWxh4ZaLlwGHmkvFE0ygwTC6SpiCYLs2n9/7suSqntdUnfBYerIHGacYobO4zPfm2O
cEUXpaunzwKHicMwOY4WhhOfvIFVRPz1DFlI4uzmUhxi31YXkRFPmaXrNpSXQ6jFPe8I4vD3SD7U
XitmLdMk9z+jmdMhjxiLVtxoFW4WgXtXxkvrUODtI4ipMUCvIyOg27TsRYmCzglVfsijfo/5j3fd
5iU8RvJKmDiDwdXGQB3fzqO0O/I/ZJuW6Un79tES/SaRJXWJ7rQcJzK2rNH4CRQq+uBeLFbUpZsY
o9xpvDx+ssg3gySg1UG+DR+HIXgnUbO+ptSJIjJg61pyOtaDZ/EwmtGXr7e7Ex7YQFsribgsD1zx
uhcD8EpphWkd4F4pJVxVu1Y0K7o3juff6nfIXYkz/UHEtFPT6jkwkkh3FZpHDcGFpfmTkApab8vr
b1UcltnBAuvKsHTs4pxBunTlknYcUthNSA5KZXvfaGjbAhl8IbCCk2g07YWIkbWuWtlhCW9nHZQM
x83UE9/w9Kk4TlryzUIgMPFa3mIejvYbSL/0RLbazC6iAR1c1URkWLP5WIm3PS89CW02gutxfdOI
yqwKDTeNTgrfyQsuS6rAeBisVqGn9wZo8t0QPmA5Uv9VfKgqXpela+exf+jBU0G26U1HxzHdUxiG
wvy5TZM5Q8PXhrBoqdZFfAoH/5YbMtZ3rViZLPGqEW6qPVHiO5nQKVZuJ3dojKsyHxBzTbe5jlEX
mzX53jUiJca/nC9cTU7+ixLbWfwnb0C2UUwaBESlRtNaIXPq2CHxEpX3tdC6TXH0Ag9ICPVyD1F6
BaArfOgyy/tZpSJU0qAYi9YCFZXiE0kUULmXtK8kjMJ3zwACR7vfro5k9uMYMdPGEb4bRmEVx8w5
YR56j4rLLVItGzWM4jZUCJNK/pWhibaiQOt9g2aYRaickBsztBxUJJ1+FPL6seuNLY+5s+9pK7qw
vfje7dqzMBoEDqNNgaibW6NJrd0ybjao32q37Vp0YmNJv/vKhAXrZ4FggQg/96mBK7uTPW9bkjfh
eaLpOvajF4bU4VCUWBfU8hBKsd8q53Xz85kJo5j/7I/18scDufdV5LErJGctsLOBiIx8pqhPVUEf
6m/4zUsgecn3rU6Ua0ok+jyLBd8o7glhjsgfRgyeQrxQjOUfeY0JxmUeSnvV+GYEPAa9ANfuV6hK
bmaLBHu7zmTPFW3NJNupDNQSxsVONEmrybOxe0K1eVV84qJUbRaFrzqsNNXuNiYA06BMy3nkVIfi
O64cmn81XWgG2ykjvsZstefSMCLFCofL9I1c2k/Zz/8KmPCVe+aLR2A1hvV5zqFecAMNyKzwA71+
dDEMIbaxPVBkmYxkI4keSeh9VDm2IipcuSLQBpYx1pngRyhIGCABuhxeGjM4IKDURDX6xhjK6M2X
hYrTKPXT/g/XSFV6MB1GUswwIG46XnTzQ9qEqYD3mprlLP2Mgp+lyBQlCjBQtT+INaMzHFbIrBPr
cUxs7mKIaPLbud5Z6v1TZed9wsiGNodX7fLXIDbUe+VHyFZEy6UgTSqFIWfmnDBR/4OFHNzBzC/l
wE330YMMzv2nllw0PAW3+83K2oIpJ2FR3ONVI6Gn3OoZEIRl/BWQtQCBeWEVmIgPWG821hUdv2ek
adW/JwHxnYlPQUwoQg3zD+uY2ULAZnCXvvDCjakbg224P4Uskp6FHRvFLvqiQI+EAobDWY+XcJoY
P4j4etTqTF1qsjR0h8mwPW4IG5d70xwtXaqucRLzqZKeCS5SY49/hXf2I3QXf249c6VqOaIiBOpr
2z25R8krljENthEziQPM58e73ZWiOFbtnTW0GwilY9soPfbmZufsAbWaVaajeayFOf8qVT10Bb2F
Hr7M6UT72DS6iDCFLWXvJFuoD2UJpevigy0lI4FD72Kis4m4WH04+tpg156nZGlM+gKg7Izv9CcX
E1U0zTGt9zw5fv3wrvU3amqqA5lBAsfRBHH9KXjdcBNZ7SMXkA6ffFSHY4S3OZZjGL/RybaHrZYi
sxxWinumK98I2N2YPXGrfy4oYyTsnhoWIBpVxWdM3yr6RonZ+ZNJ/XyawYd/VD90SeZ66esiJMxw
GM9HZTpSdAQIhL3wPsv9pt+PUrDpkxigOruTFAm0aFMTFOk0RXeqmJiVcnFeq2XGKZMJDV16dKYj
ku9T5qlJ6vJZLRseJw/eweaGIhft4Dhu94eoqQW975FTaXnoNhpIRj+p39++8Q9mxPB3S76kh+sc
NxTEvzX1vkSFH839QhhbN8GYrcDFpycxDSj9VPhQgwMgVwfXPiQQhjxrfGqi9tqb8LFyV+lF8p8e
wGZHgj5e7EdwEJYjIiM3fE7UklgogNFs5d2LA16w+tq7211+r4qpFQ/huM6PjF6lFtzma5TmaRxh
+ZAUc3sisRjXCKVWPMd91QEaq8tMmAbPWZT8r1lHtFlxHd7iKnmFqin4XO1LVzPKJ7KWd61lID4/
j33TI1Di0jddCNeGOrIN65yvFwdOuPOrs6sG0FWaiMwdG6ZqYrdOMQUDvflFpUCujcB+SQPhMtaH
yETPx6TBEHX/l7BkJOkLX9SVv06Pd1rIGg3KWJwTIvZCVA9TQRTrzfpPY0XOpoWYOsSBxSMg0SOi
OtY5lELWnN5KD2HHrjjJ1JmTEGmWUPR0trbZgLRDa2vqVQ23VvUO+pejE+WhrfLl2JzoOHUMNkFX
knr3rQEu60FScVxQpTzPNnY9RSh98cVPqpfxXuO02hNVZOUH4gjjYmeNj5kXbLNZQU3t1orlD8H1
PmYCfvyGUSdZXz0GCrpzReHcdkyq9Au/EfEqwN37f7paAGJ3z35q+N8ciQptTQOJghsSzhrgxj2H
Jx7+S6P2Y+d5mB6XK4MxuOEUC/ZhUwR01Eph9UifjtVGd5wvXzLlQRETTdWgMEh9F17PF+XAge7L
q7ckXaksTsYu6kd3dd27E8OadDQbrzijF8cQu9R2M2aRJVjg9ppv54Ypi7wTWvNZN3HPhxm08yuW
3wMaXR2SMRI+UbcZONDFEh/1EqFvld094FzzQSf6bwhX0kfZWCJNQ2FYshOGlMGb61VLVBllnEdv
YCbHXK07YPR19R2/D8Egt0UUjjHyw+342cXxl9zwyV2MyR/tr/n5M3CsWXyR0J8tb1RkUQhhXL/p
oVuC/2P2iKWWZb8npUAz6q4di9uenpe03+o6MdIz1cZFFLTrh0oUGqLOLpU0cEaB7v70w76tpa1F
o2wiv/iMuDaWuYCXqAGwqQNxX/u04mqBzVPAml4QNNIIP9P6jVFH7covdZbddlyehp70safTVhzk
qwh/c+qbjryIiV6TGlfcSEI+PiO5E46kGF7wDGppOHnxIoC0i7sGJhsxh1bd2tQpv0DEELd2/w27
mkdq3JMekc6+dRhFdPMG4A3bVs7yhM56wiM4IqGpIlt1ARnVAExymosKYHn5Dshp1rJJ1YHmi5BQ
L0Uj5WONXycd87Nwr43MBY2QzECrz0lv8xuhosgLjoocJpNOxoS9RPRK+kc0z0pOQ/ykOughS2Ky
1Xxg2VZP1NM8XbrXlvNZlJH4++7YUOPUGh3p4ULi3pb/UHHeFLZSCmygE5ikD9X7EQgyVHDEvlsE
G3RbIhAu45/uNn82dp9aKNQ3PAFLS6qdEoJGmZOImbJ2GvBkvrrWpR2wsm5JFMF6BOJ8QXK6DkCr
wxw1Ju19FvC5p5GAq3D/A5X90EDppXXXWf2hHUx4c9PZuozpzRNMuFtai2NIbeFt7gu6W2KmsP81
rnysYEqzVuyVsKzdEilEumRdBIBNRYDo9kUn4dcpOc5W+2QMX1ZCzfQi1E2hONvElxnyM42Zye3S
8l7svfVLwst3AqdDhrHPJBnhDWnjDUmfYbe6Chn7I0Wg1P2rD9flZoCAVAyPBlFXCwXOVuNzd8jS
Ws07Sa2o0RTwHS+bE+6qDmQGRm//hacT3MHgJyDGM1QrOsdHDmTmGmMiSsuSkDNmfBZGwqHxM+6Q
31DjBpNkSWO/zmGtLN1Y+U/9aXZ4Fk1Sk8yFh0VkFKl3vW5ZSQnlcg2kuwMK+yYKbSj3CLNqat6r
54fE/96nubFgB8xaMDLQkQo0dCt4i9I6BnjO3cDYSe3xbE1m8+EwszgbybC5+f0d/JXAtHRaIBPC
7yduYtX/Is6LSrk81L4+WcrJBe/esV3rvAdyNhLVmAnw5hDjabFwlELIhsfn5M3Vu1Wi63AgUH+5
/rR7dLBTqJPa25B4FC5gxm/862VusVZUMETu/O+gXkYskZsT6ys3Q0Wpw/YS8PNUQvpOM41qLp/E
QDJvCLPKrAZjjxCY/4GZnLN2PXfLBtV8th8bbEN8JKTfO/NRRUQUGkHE4pnFpUR7iUIc4ssv+Zj+
ztuBh89PWjnuOG37fRSB4qRt43L6hImLVTugroNosv+2lG5XcLhZ4JDAweavIaWLoNvDKXe5u1p8
6ighU4VLF608cOYEWqDT3oZut/WtgA9TOQQFjZTyCBFe9xSnDoCox38xNTpCSciCAZm+ZfAt/6S1
a/MYJ1N2vkslq5nxDOGw6dDsHaxDhO1NzjtsECaQES2pIIaBmdql7y/+9No6libN2Qvc1Go0SobC
y5Z4SKaUhML4WhU83RZzeNXRruhHwDz3Igrnkdr7ObfP0Zbt0mNRPxn87Dl6AOLUcSWUa6Oa9mDz
2PQ0udDVVKS+z9LkYvqK04wAb16rZhB3B0iuqiDe+0HZUKZhdhlJznXj4SFvqGiJSbiVBAUyHymA
Ey/FdeGIhU/S8fHhJ38lv1/ZZOXc5BlSNe/NcDzQV6mJW5xCrFn8wAsjvbsoOnJRB8L9bnxPvyEm
ArNHfJ8r+0YIUvswjYcha1AgUb6dTR5MaiE40uE6r5wQAS2M5ooQxvePp6roZ/eCaAz/ntmZB2sh
pcScNp25FgVkt20rp6bjd330AXWhbWGHohCnxWMyc1w/fk5zNefkNcsaNWrS6a8xTjsoguT2sUPj
o5dC0cazy0jBghwWDC1y4fLy6M9mwRBYcDfNCbOLVMinFpM6ynELAVEEoKKF0k6perCn1qjHgxeI
UaXLAj/+0R+IvexUQMpKb1SpfV2F/idfXkO3D2PDXr6fMQ9l7Ficwc0t/0nWpEo9wsirYiLU5dI3
uhfiTrePbK/DwE2oYvMO+fpISavV7ked/n4L5F9Hl9OZP/YsXCzunK4X91nXrEA4Wf/cZ2pvwtKA
wfGXwjn0SB+6UlVka05rzjHZvInwGjuq2wYVMaCxvQvgRCsuf3p4FBMgRhxJzSZPkoIaBI2P6dUp
6gsZcXoEOqlwfh0XyyTFX6gpqukpOzdsTT9iYIoTDN738n/zhL2AHlPdOrdv/0ilPFmTrKTX0GDM
7RrXDtY8n71V+hSxLtszc+bj3+m6q+s59cy1zgZoVBY9naXDyazDqlJMHKYbuC1y59+d7B77ra8k
YiqWndCe9samt88yNrFPempILcF1PIYLZ3ak/kz/weN4T5As6EQzxHDJPjyLeU46mQs7ynekjEYH
4vSuT+zxsVGmpPlw+8o7kNvMCQ2mWXrilil4O7G/xsqC3NqwhkwFfc8qWnKutZJqad/fmwQ3R0bI
faRe1yxXRrUxYHC9TiUm6S6ZhO3yr91Ie3VP65tdcrutgbzPHeEr+1m6XY6sdsVaNtJcbAnatFNV
LiVO5GH+/szLcUPcQr4lQ1+nIzhM7Uv73RzR1u4vsQ4qDOLaiHB2k5QjZMnvCE0Qf0IYh/ADnXzH
OYTYcvCTHfXroRFjLc/ULMnIKq8KD2k9LWJBPb2ynBdE6dxTLrgWi5E9e0mYmHB5M/g3BsVlz3Hi
LVZXitdETiBEstLZ2umtCIPRaUqk19g+/iQ9Qc18nAXokWW3ro0nfNp/KMyTZqhWFtlZXKq6+QPf
PNQG6DStwBP/ybyFmt5XAhP3G4rta+i6wapXUs/n/kPVna3GOFA+z3aMyIWocqA6ciPdzSSxZF+V
hnEtXt77Gi2MZ+XyVZSh5dcg2o1LCFyi66MQ31DJshVnUrBfSwqT0MFDc4Swb7Zxe0cOeukbtfLK
Ily9rvPSw7EjmDFuVnPcoz6Ca2lIgwxz2E3AFD+H1ckImQmbOFx0iM11FHuFtrFQau0Ey09jp4Jk
KEoQXWB3+S9eD4a2i0nOW4SUIJlxqDY3NjnjOWllpbzdHw+IHD+1qbIcOZaAWLqT26c5dvpYaVND
x4Jqb+pN16V12z+xTDeflyOU5gBH8dvzFziW9W/I0rFwO2dWVsIZufsZ70tE0Wxia4Xj+DPMZO+J
NBEUcDJqN52xGXSbE9TNi+XmSMyCJiAHb3BIm7VpYzYylOfWe25V0zh50DnfeVhLjRxV2D0Cf4DR
p4UlV/zzbKB3AhuKWgiQ8IS5VX/guqlc1liOkHpn0K9UHFikEK4JYJ5z8rYDZ4+WhLnK7MAUJ5En
TOaEhrDWalQBeUc2Oj5BlOnZrC8N+2CRUA7WUTLqGsjfP6PJREuxf+eNcX1TnvLqvaRayZNIAHw8
zcoYzSg29ztqhCTunJMJDOiHFtqVQMbDCW/KouHhLuucBqjpqpR53HVga5kzbT2cByr3sK7Yb/Su
SB/01+valjfnTy+4gv7fo5QuKMLLFsrzSCRk7lZXghLmQP19+ut9qZpHZNmyD3stNMji86uNnNx/
oQwWm43Czu+B5AP2zflP5mPVP4IlO0KLoinnN0KlcrPY8UfMJYMT302JKqqFDN5eyltt/LKJhksE
xwPrQX/Q2hXaFfQPJs9Q7Ch+tOPQVr6/8oP5w8X/RQVIZpkgdB1DMfiJBVARw2zUYyrT3P4/4aAn
LaE8NLFabPDTRKV01cd2V3v+Vj39uNjsX/p0YPo4r0N+Oe813k5xXtTDs/uzfFL2WjH5bYeVP+ub
opnE4HmhZ6mxFke4VBrtK6BpXdQSicjkFWFEmGXctQaIU5XLFdotaSd5l/Fc9BOGLob9hZ2ZM8F1
CTgaNIUzkvfDydDwPbcd03N9IiSJM+J836msUeevIpbDGr+LlEoDIOoHN0JcPuHvFkGokHu/bC4G
b1icebJLjllPoSTYQxJIW9Aob3g21Tg5bdCTRCYa4boGWTh+VdzyhhmOxp7141+WuNnxtr3jd/oE
zbqPW6E6kCgO9iy+QEXPl3AguFd88IHeC+80hynUmvoFJqgbMb+YtnQo9W6oADIaByLyD5IaIPyV
Dw0Wx8rX2UxJk06r9ZIiQGcP8YhMBoHNltzw4bAQ/IEtzohw3XAZTqb/vEsWQIPpB9P7H2Al1Cgs
0Zme4Rtoh26QYTzmLw9ojGOwSGy34InIuIj5hGE/FnAcXyqSqCQAWQRR/vIbHKblf+s3c+49xKz4
VObpOEoNO0SJpcXsDHL5Qe/CVYt9lNVqnp1ESw5GCXulOiAiE0/zZRhVSRcSCU2Tnl8nsFMcdVpY
5xkCvj+AddkiQenHZl4JgqfjBNKeTb1gZ9XLEmlSDBmQYtx3GMyD8Ww4FpOq55pIjXzVP+h+XaEX
fhtNl/vhdZjsJ9vm7u9uW0TugnwlnIxT8g2wo8VqvGuKklxqAPoduPr6NaptvJGIvB0cd6i3rHdf
RhXPsju5S5f2PgxixlbLPu8Z74jwfnIpKQw0tb+WdE/KA4vgKYhLZB2BaZvszliFPfDFRqBT69PV
ZdHlrHzMrMrR32ZKU0ada5wJZpzR3G3kNyn9tbffCag2XCyWb1vq19qeEe9TXBN/kwXycT53A1hZ
gb2chesh/zkhMe/ydOeiObHdbiCnUgjO8kZyDtd0FlULHRdH9dTTj1cS0Xi60lIy4VTCn5jSmeP3
AtQDP9X4guhCPxj2I3jjzWHnjvZnAbFWlC6UPYB8MacM+RemyDLt13aB5t5bbJoVhlVHqO44HY8U
Szb5B/KICBzmquJNrr2imJAsyRif3UBiwmvHxesW4i+XPzs9NaQeV55O6XL8UZ1NlfylcFaHdwmy
vx/Gc3CfZNGAWvXmo4B5D3Grg1cn+cn+WqT0gr/aytlNKICFOW3asuqFD1vgApws84xIifb3TXcK
rBHph0203ZY6J5edyr+dd9t9kwY1wpmS5YAwwAcfZ9kf2abND4uHQoMB7fGYW6ygzN792Y+G+5m9
3d5DH2/mw5+tGtNnqXp0lUej8HvZXuH+69canIw4+JEaZqdE74KL1EhLQEDdNOEr9UOXrycI9Xoa
ec3k6ltGcicdAkTGwOoRaYkfFNMOWJfzc5m13/NeGgBelDIg9/Y0lwyMCLev0oUQLD5MD2JNe2UC
eHrRWK8Z3EfQj6QabPjWbGDs1HUhMLpbDh85NBAM7Lt2kKeO68LcPJeXBuDZUW8JXYK9WFwERuCS
BtRnzxnPu/zfx3uMjq9gcSEe1MGChIPS1ChKGC44wjZXNfscK00izunZJLwTumr7xJTdha1tMS+y
pZCn1RBCsAQyZbhubGLvy7MQXpWDxemJ+rhGdaNPZJTxwIt5L/LgNoWwXoamJv2NP8HC/7K65T+m
jGxhiV2whjwmI4BMef9CSS5oDI0YBMvqjzgTqF92UnfhzBakt9mlU+bB6KP2/wbJmbTKQAMaRM+O
YOi306R5pwmla3g8EJ9gfsnkCx1D/5DJJTSi4OwxnXmKRDFw4l874fnzZT1HGfUYEgusmpRQuFPo
ZHZNN8eSymBAycCh9lF7v2+zH6P52wmB3L3/QwiEuIMeqCTow5G2rxjwb0Mkt5txcjtKfSWa/xRT
X9lfk8XV/s/iZ9rtYQaAuqSShBll5Ri6FxYjhKDtOJxMx81wv/cVMsRVjh4vV7ex++fuFXPhnLs1
G8U5FxGLe3/Qd/SipbPc2OWn6P7EME3qmkLszmcBFJZfdLV0RocxgnySxMM+mQb01DKh59HcRzhr
JlUW5QJvqcRropFsn1RM9XTLG9EcxfNCTGsUAiee+EdD1ThQL6lc1KFm8DioL103Tb1ymAXBpFvs
ura0OJNVBd5GaOOBQl/wL4QYWfCHj96krqehAgaDAYfRwDOReVXuzBQA0ufJKrrbhW8NbZEvh2eS
PF9zSxq2Itt9pZ4zciirYQTyE4ufJIIGS5Jd739whWGBXOv3KhM6JDOVAf/mEPskpgV6N4OA13pk
nQ3jRo99NWrTM7Mzn9TjYCqOrdWL7MKsVxcC9VNGWvEw0+V33tUTTdr9nDSA9pkcd2dM/FlCVNEc
97Qsfxh4x8oAUZ8brwIHVl/cqIIN26Ek2kzJZiRHjSAEAioQ7hJASXkat+Q8kkjL7J+t2M9qekLr
lqaZIknek5wS6CJvBQowBdWfUdBG4PoUeOkTHxJuWNazZTBBnS67x4VK6npqgTZS9ZuHajO7VQ9n
vjMAPGACrf/1uGkWVjs44/ewK7oHzWlLGdinzWYt3+689otdorq+OPoDIiK0o6LQaUoEW0fu9N/K
lXJci8TSI47KHvEFq9C18t5XSGW/NZ0u1IWhO3sNd+7JiF83QzDvwuwptq8KuZslv1cbzM0HYFrD
Za/5JvGo2Mdmqu5wPvTHbmfnYMQNd0qrt/PRrPob4+xdZBTkqHWVAB7nfdqhyS0VJE4sIUYlXxPo
7nal/jcGeF5cHtbdm22DmCJABg15EWR/mptSUtd8GMdqk6GBWgg3OEySlXWf/23z2s9gbi+nQWGh
Nc9ItTaH6vm2qF46VlWCjVw1PQii9eNZEl3Ry0svlNFaH6QeD5Lt316Fs8sT2N4tyI48v2vP7Rr4
kntANETkb3LNFONtYAQarXFVv8u2WyG1mlXu58x4xuue8yp1VuPGcBpbKWMkWkexqTAipX5ZP/4F
FKm1jo3vQB1CwDj87w5lAyrbOQv+dK/xPxPAZcS/hpsLG6Zn4VyFuR4JVKeAhe2QMBTi8MBpKUWp
jr+bZ+WrwN6L6fvYZEIm1OM57u8Itu69OWZXLN4gVuKanlPJstbqYzvAf2JLiwBgDmZEjm7dLFmH
tnNx2qoF4rslI03F0awn5TWirSrU7LSgHsZMYeSkJK9kXYOJPBHvkW513eywAAV4NF2iwZg22wHV
fwUA7tQpyATgMca9B8hlrXUKQpkk310Apjd/G/xfNrAHnJx29OYIS/76hHS++RfhGURAxVfyu3pa
4HFXAzlt9dldcom3oOJ9DvZYD7gy5H5ZX8Ouyy6+c07H0mnDLzMJjkkWwhdNNNcpnWZqVwR2hl3i
c3nmtU31a3hOoDL0UXxo1tswx8cCwceFdJaWOTXy/61Qz1tqXtnkCDj+AbMxjBkviGmuXKfnLd2V
HIX8dAGTTukuXk4C3PFMUtZLNCiHV4MIFd7gok2B61tfcJ3a0LP1+cGUkrzj/xpznyzj3gQZpqkR
4OWveGi3w0aToZKUPyIjKhdKlzuN4Zb9Q0HsYQmCMS7tUpRsNSkKqkO+Vb0CJocYUx3BpOORCDx5
ip7f3qU60LtjQMkdfNLli46vv5xB1nX0PNaro5pRSniMhnEs0wsrlUck60Md4ISzKgWo5qucBf8K
1z2Fno6Z3obtqmhbs5qMnMOcnt0WwEBU/FiySsQSbufyap4M0i4z57aT6UazkOBb6eYYYIJM0UMC
/3ysU2lLdtOuKDdeESbzmp1xKx8lfWZkCb0YJ8p2rmKyObnc+N0HnzGcEccf54f5lE8myh0h38jH
YvaafmLfWG7UXw6AtQ2QWg4CZts65/GpLC4/jHea+zis6rh7fIU1o4FZfUYxJEktcb3G5vSXjvWe
EUSQLVrFJOpZu7Pj496wGWR070oTTgbf1MEkMyXX2grqudd6Cx3ZbneygLiTd0ln6tSUDySwlX3i
RQMzOBG1nyqSGrdbNz3GaUPkcTdBdjzNZTKSrfbN8uI+aGKqOX+qp4eZJSRYwJecSMFCrmELpj7A
alyBtddclVPCLuMlPuXxALPd0OGv6XUlUwfLPckChONgfHzmzgVmEz8ystI37fOLQk17ekYoTBCq
lVpeRupUopbBFjKKMzMFKfFjSqi4DDcq1N8pYHXxxEr7OGBV8wOXpOOL+fuwk49cXydI9MxcC1Sg
xAjQDqSMq2ARoHdNo9oBGeFd8tWRWLdFDjTWZ3Jk7H301NuycNwILlbv86RhjEhWsJKS95MChHen
HL9qHYeiv6ux8GzNEDcjwJGIwwePHohRAjiWHVT3kFpTmg3D3Ye4AlXhW/dZhDqWXXw0jZ8/W04E
oTFlj15H/ARTTstsDn/nScIW9hMfSkwbRpBTUjkySLBZn0uZqF1Lj+rTtzFiQ9lOvCYouVdprqIc
9SkvmGGER2/KMhxhmxVZoBoY/QFOgWw/p4wd0rK8HVUckLLEUZVB7uzm58jK1QSdnaSWyHTDYQe2
Fuuj7EFYswdVS5qy18LuwscWG/kuf4EMUqRnIPtfF4tXlEMtgV71U0W8oVTF/55G0qqssdChq7im
vAuwSjbDjmQgsWH/z+5Jtb5SM7fMNtcV/pCFY2OirUH//wLiQKoMcCu3ayQwgU5b+uMuljYJoYmh
ndzeq4De73B0zE/1jIKLH3GUxoREpQNKCCYjK5aD4S0FaN9m6kuA3xeh2EhLbxHv5XBTqXU4V3qq
+d648FQsDxCqCGRJZmMNF5uwxZFsyhHhxUsBYRNhAzk3wXFS8pU5pAqyH8EStibFoh0sgRRFAbM1
6JwYBbhTIECEyKWi20LhU7NMcqbef2QKLketpD206C3Rp6mulZhFYjmPLL/CAqIrOr2ZjOsiWRqn
wrgQ8vE2EYzRRlKQZVSr5P61leF5TQUqDTMlY4CsN9Rw3wd/aXRfrx0W3jUC7oUif/LNBMaons+y
JAunzD9Q7SOSfu5oXO2LT5BMRV+cqjSAEnRM5bTfSuKPH7ydYFO7NcAQg2ADoZ55cuhC3xRu//fa
NSQQy806kddWY27+M+zztO392kaDXuRubOgJjRcc4qpIyNY/CPqrQ+NBW3bVN99Yyx7Les2vFf8M
5V6nn5CrtyH6KjE9lFQ6gL2Pr2AU8kENhHA3Lf1VG+88gxyTfGHEzZvfe6AEM84DQ7dzxf3IHEjQ
hsdmM97lTX6ssZxw6pOVkvkyXDLeFzjLP+XNRiVgIjTjqnK8DkDXGJa5Qyqg5zpHc+0SQpAgQGwd
DDnE8iU4LB2k+06YK3tUE0TPR+fr2CFMZtXhx31TD8uTWu1Wsl4epRNk6G+83g9jUTkf7d6H6/7w
3TtysK82GeYRsvM1zmvuKeGu0/hOw4PUuKoEW9JtFgxHkFY4gCzbvJj7mn+/l0eyskCTtGn9U+f3
7Y5TslbgBObrBcdGNmzeVK1TJdENTBvXqrUEMsC3uPg/rl/pjyIjgCwwWxJzLhwEWQmPJzIAZUSr
IxkePrEVtcYzQ4j1nEJuanpXe1hqhBjnbllrSD6hteyQ4BhTOtw6tInNQFLjgXice1aR4GNI3h2D
4dgSXiRaQcToWuGsbRrutZHqqAGf+1lS/BdCPtlJ/89fvaEvr+6DIW+ewFy0heHKkxigj5m4C+n9
TeUZdFGRI/GCYXbcnU4qRujsEwi6xwqAZWtXM7nkZE0Hs6vdyJCTXoSCvDSe/3fQjJ7ISA++Phef
LmZQ4woycpRY+Z4xVzvoQiI3qDg224mIOe/8NlikPGUOdTpAosC7fIC+jjqjj2m10DIKmLv6Hua3
O48N/INsFDeEKOAGGJ1991ppNqcjqSRkxZbexkS7DmJh8AuAhDTSeY2wMXwLde8BPU05yU6r9MxU
VuMa4ayQOzbR8hs90qWNfXwrghat7yPPKmucXky1a+no8kfHsIMy8TmLvrfeQMatyJfCs94UxdmP
HpLcgIyeZMkWff9I3SQ7aA97pHlSuxTIQoecDWlx3lL1CDdlwrHgyFS6UJWNQo534LEz4vxAwTAk
grpmd533t3YmNE9ym/CYHQFFJL3DkB41Z40hE0Lrq4srjhPluW5J6IAyVFCH1LsXWv7TczKhnkm5
BGfXXa0DtWfOSsT/z8J4fF7plKKErhGWUSVkE72qWkgR7GbFOGc0K5n5x0YqiF1+BetIIQ3/Qwe4
ERHo/jSc51LnJAjhC02jRBrUXijpzcbmNez2WLHBBxuhE/kNSDmzF9c4qb+UqS/RDuuVJZ0BAVic
JtU2D1EWi3SLF0MJb0czX6TA+bOkpxtNCNMr6V4qpKZJ7rgZmut2WEhTVekxQtVSq3LPUUQPavOC
JwzjL7qa9N/z6XuIwXERepTlksFWNureox5xt///A3BAT9vgxm0ws912xu0YHjQQIz60WA8KTGcq
geyz343viO2mBaL3pyWEY2k84ttwlMguJcJk2XL72xy5RkoZ3H+y+bmT4C3bYjwrrzgIdgKUJhLp
Ee+PKtFT7J+ovKedfYVFmUI8gfeqZbPHB8IqcxH5CPIKg1CvlbPHOhImUH6Jv/mqfig8CQ3z1eW7
ofZDyR5kpFmiIDAwn9lShJfy7dtVGOgn7geCKxk5jNxKV3eK53WPH8JCbhCFmRm1iySDli7svNO4
zNVw4yWjkBwY8IL07QKP1+6foSDgTdWEgmU41/+BursW5ZW3AnBR65GGTq8qSYjIcyMokDHXXmSw
c7bjTQzQz2NsTitZWO1W3lig5bIZXQjDkMP/mk4MjBNIy4Nl5XWsJbfADjL+RIAqwg4IrsXn1CRc
8wbv6Gt2Kq0ssIz2oO8vO0sVvwaXziXygUgjA9/oSVf0DHRWB/aoSJTSJ2aSpBzY8xa69Fi5C5B/
67KgPhH6RyfhK31sb1u5R3ePJwo8HRia7h4W9yYgD1k70ny0BxsynEqM+okkirijygt7EpqZ5JG7
4vE2/mdBjVScK8Rczt1wZydcwKZ6NVSdM2s981ErAEgwSsQpBRdxhIKa3vD9sgmfU8qXHvog3reo
sVUIX+91cmTevASNaSFcCumk5/H5LBYB+fwVxMKVKSjrTcmpQfq04o370cb0CxRkls7UTvAS4g2L
EdrQnMFG2ur2UUYcr86bQVnUoJ+2KwVzzr977hrMXZDDdtASWQ1sASHyDAzZwbzmUVimzQSZrVZw
WshnpOTyvz77Vl5ikk/bFf0CNqauxcw/NFlb80ZY4JzYGax3dTb8VxNqMTE4ds08IBI/CYN2Pbqj
+whSmq6jJG4IjcEYFIEq87l1AIbdgTVlf9jF8c5QH/KIVAYGw1C5HMFr3FXaiCLWB1NXkEOsK9mI
9PmPEkNL/gL/te5i4qd0vvVkvUUXTVTYqCenneNheziCjzaOHStxnvHfIgfT42QnRrE3Oka/VEvk
4HmL1fjal/EtIDACfbP8x+2ODNhGtUvKVGaKafzov5K00wISZDX+jUkbKaAw8ObM9m2NtGWBEOsI
RhkSw67ZnogvI0Ju6Ob5k0c6DI9cvn8JD0mmBVzmuy66fGUGhqwCRy4inyr3UiWwC2kd/HDAzMV/
3iTeFiXQj3DcV7UABY2uVGOGbIPoNw7ps2MOjQVfbBWIE2rYVNmpMzMJVOmIkYG26iHovp3u5YAI
m06kieRF9BCEnXv6Z8Uq+C3YIU8Hl967/ku06xepGJWg3MLo/pOX8ydohPJZEZECIV1xupZQZpd+
9y3v1UqsqyRa8vmwStAfGUYJr/BD5oDY3vc2OEutiQS3NcYd7QRr6DyGrkrEkpA+Vj8VFOL02vk2
Q/K8BbcPCMDvk1KZkN0tdedmfMMBfvoktnNyvmmKyxKFBK6oKmoq7IJbeJKhJXeJkjfCc9z7rdvy
z0DmuGC7IYnlnhwadVehRvykTRzCbNTtk5WWPJdLcAn7kQkmtXwFBRuX+67yfM62d1QwJmgEM0KI
raWn5B8kDePwSKLMkE5su7XDqkCa82z+Pqrbv7vBqbbDrH3pW3c1BgW5iPxa34djLr+o//CobTVQ
bGOjkdd4SHPm+HjlHPhPXVhi32irerKvmL7CtiOJrbVMbQyDzl0P7ls3ebzMNna5gIv1d5+ndLlG
h6UPVKyEGPTwt8xULdN9ty21p1KhYFdNdoQKNqFh6sAgWBQz0MSotIcUR+Pkx9gdFtYJ59bXlAhe
iNO6ciXBO48py2ECf35m6Q/vvIjLHRhBOevgcXSt5dCnVKpbe9NEpfleb81IlpIlCkpXxZ6J7uZp
w3575mVckPqxDvQQS7OGlTJsNWPNsDOUkNMfk1QNSQl5EzFKMwc4oRgB+0tUpc3lQsLiBQVu+Tod
arjE90GNyqA1Y/6jeStLvHJhZJitC6zihfrysCXRuLWHFDaMklE5LrzpAexx3eIvE/i7p6odQD1d
BoGfBy1/gF3qt17Ns+stmuy5qTzCnqv65B7QEkZeGBtnpxGuL6QCxqU3VasbSxRIeHshJTUox7ON
Q44n1MviY/ix0xQAMnhAPiqmZpksbN6F4MNOej7i4yduq7m0hbItEV5+kuWMb5/kNCBipcydPpJZ
HyRDnrsbQ+bXGoVlP5lFbQPGh4b/24CS+TP+eQjaNB3SvMLonrvtMl8QtGU1J0QankAuHh0LAG4O
MEOpaOFBLk0MbYaA1aHmXh0l7mHWzoyr5FKAv8f1ybfuPla21v1o304+ottFdv6LF2hVYs/N89me
Dzlyf/Z/0JVZbxOxp6L3C/iMTOPejv+UHYb/+5t5mu7FJVKvNAvflPjGwwZmOy9xfzqJ+NPi7VDA
IhPy0vCbkwqeVuqjB1lvkKRIqoLAyKebsF5Var9N/DpzeHfGUILV8T10EXX/yFeS15SZ9LRonXpc
vP+Bvov36YbuzHpqFJ98dMKN2+GeyJuocSgYYlUPiZGzm5mNlt2n7UjzknuVwWskukw09C65M+ZK
preHUbFNSVfMhLw/vOCwia+d+GLopsRgzRAiUS43Swe6+2zl/XFq7JHhZIPF/UYahYXT/mijcdq6
M2ueA8g7crR97ELCQhDAN9LLBc4xvY3VMOfVdgMupUGPlizs3euItRJfKpJzb8mAG3jfI1pauvPe
5fr3N4Z43x2S40ioLrk5SOD/s4QiC/ORHvDCL/A61YPIwMI59gRHEusBvYzI+eVDEKTcsfM/6HZn
GlJY8gLy3Us0NShi9TgXVqxASPqo+wOAQTxF8rq2S1GNODcuJRG78Eh1gsoi2oJKGuFoVPLCdxhv
UKjirdJ5DoJD3petz6oZDxYTtwZYRper8doxE1ouZbwfqyg6K4MG7U4qUghepm4PrpvN9KWsTalK
lWVR2/bq/Ds5/ng/Lg17kUpqDLDgK1xs0xDO3stGvE+QTCpp0D6HtC88v1xs4dCKJooZKjBmE2At
0SdDdO+sy7onWiWsUU0aTiz1iPC9VmvJi2V5gGY2PAsRXd8WiBevqIDGM5Y7aEm0PjYn/bGCSusO
4r8RRmFskqaYdGwJ3/A0eWdHkriaR8CAS4n6L+ZwjWkUfCWN1/VEUS0X4rZATzmWqtOtGhnc0dxm
/TIsrBJWwLh/XDXigMuukS/Au9y98DFGg64pknPYSQ4FejpRz/N15FEiPAZzT19luvQ6eDWbEQR+
3Gs8CxXQwlx06r5bxntZgNZS1jOtsp4iPDt5c94p5K+zVvU4lDX6Bh4FoxrxMg+S/ugsgff4Cm6E
bmhuoaBC4QbZz7wtfT7ICSL1GePjYcBsKhzM5DuwZOw0bWNTXH5Vx+EVSm6beLA2DOw4NQ1loyRy
9I4sw2N4ohiUl7B0PpR3sj0dZSDJbZbPd4k2oZd68eVtwVsCEsyJgZMgAeOcJhoX7gN18alBh5Y/
IsJCIdH/IuUeWyNOlQxgd6zbL819MOE94s6t6+fAa1lyFfAlSzGiWRtq0XwSm83C2jMgd9Utscsi
BhFeWPrY/6AczT0p6kD93pe/8nznQZT30pcxWDtGbPBaC03Qz3F7da9Xy3SIbz2/lwTLhCtIbmEw
nx5baVJ7bx16VWiWVdPko7coie6SgxbjWP6y1PK/j89YHW67xMy5iex3DmcK+qZ+MLOoJu8CRuGy
uZMVs/ISWP9LVwGoCFs1vpt0+PvEjj442/VftMUkD1GZ4d9FxtMLMknUkgJCVJK36Wjcasjn7HuX
XXs47MiSYMnGknYWEY1jaigp+Ri1BUxPGSpyIVefXMUoKIJ8+SX7p3NqnmSxsZHlpkCc1sbffM37
/1jNe2fKtJ4uaKfHYhIruJmxlXI0wCgxBmxKzVUhDTM9EpPSFz5BO5CCFnzN6A0ogAoOHa2ZTpv3
q2+BUVNp/zqTyVyh9m3BZBFc+5EyGgEfU2qGx+/wSudCQU6Cz5r7tsWzvylf5iVysL+h/jGsbjO8
WkksQfCs/mlK/qDW62k/M8odFIqZl8wcMtIkgjWpJuIL8GpLI/qDOCx61D7Dn/EMx00ydy0ANVyO
a7Qj8HAu3Lnb9sqlnd+aQEUFvk66K0SCJeiO0rrdgpWRqrl3gHE++B9RypxQBFO6Ic45fHac7MPR
/IONnyv//6i7KTowB62Jx/foUsaXgg+ALiF3yeZC3lyh7IIIXZ0UaQVuK5KdnrkgKj3ejLPGpG2t
InG3tnNYQ18ctlwXKb78H1vA46vzy65C+YIQlIwMeJdjxN8SLwaUQBOSsTRBL4h1u1mf1q4iY+2B
kOENMwIiMXz/BxlFMYFQiAPZ9szowFWUdmHOY9oQi3pPGsH11mnBCvBW8iPqMPnhFeGpnAU7PdqT
y6bjL/i0XiexrD3zhnFqTNjPTZptAvayIuPkF2Wfj7zTUETO42Y1bRrNvOjQfFMXUlLvcWnD8KQ7
m+0AYjG3mZs7hL2z5kah1hLG84j7GRgqQe+Fks/vTkXnnPrkG+XsgIpCTkGVWJAlKNiUbTFN7sUk
LwvksMUWio7KD0CzkR2uBhRyPA7gSfYQb6HHQVGWZee3g83NDkmbKMJYXvwOCVaYYxD54922Z4Rq
o/67Vg45CL05PWXcUO2sjT4W8w8C7VhqV+GLP8YI6qFcLjtCFWxXo+iebddC7jeYKAA2LYCoefeF
q3qNz/i0iiAzGGNtu59vEJ6UdTYM5445iChxOwUwNlaw2ejsvmvMgPBA1xyQMySCb8ChqaVYJMPe
4K9Fyhk4cv8wNe3gaUl7XLGmUUo358hDx6TAxy5M5UIFe/0taRTqIOix1pMYM/+JYypln3X6v2vb
QOQSlqWnCvJBrkEt/a4Y0zfh/65Wfk28VsXdh05pwn5SEUR9wrgix1uoxZYoyTjmKjoHReupZ6mF
h4za9KWCVfpQKfISsRz3vFOwbeEKlDbKJirpAqf7dRWEp7DiMoXSMj3R627JGRjGqCDH/2Dhu0oF
ylc7LPyBBObqahI4FvgF+6a+wf+Tl7JXhUXYlHbl3nZygfILv88UKr+UhIGUTBjTeJy0GIZhCHlv
8/OGmcAS5tfiTS4MNI5Pt6u16Cs6n8sGn/LFRmUVIHK+xXG5KUoGprYNbY+bVIw6BM7zbmT7mzWF
81iCR4XqKYeKw6Jtpb9KMcpl0usgFkjxfnIANgtw0KKN9UzaNyICeOGVLa/2RZ298pcmDWIlKu/o
6ls0TjlT6f0+ddZcTZIVFiHaRvmrhWksBn9clMQkPoG1qw4ZQqgnjFxq61IKMTrIDJGVKesj4JRV
BuDfyEluLzJczS21pLSmjZgTj5MP6vfY1rZiKaVI6kapJty+ziE5D2KGxuekk95D2GGCU/bDEaSC
ZFGcjzC/XNVvYf7JMPkkGO4Bm33A2tY+ab3CIGmId/ZPoeptSupkeuXdLyIC/QzlK72wl6LIPtrv
/eImFyB9rCZs/pnvdmRTvSyoDtkmU9P1aaQrrfXbN8xXfYZ57Jisnglw+Os0fZ2KECK86K+N8jHI
63BN1pnIrBAuHxXWQX1sE5ntR84Hr4RPYJI8UfGRfUPoLh/ENDzcAsCPYW9JZSHGsOqTI2Kdx6Y/
BoIRanWlL0AYoPq1NOuhOD7hY0RZ76p+cqSUfpcbzfhZEWKvLGzYzYaFzFq474B9MAJvF2gBa2YZ
Yj8R32PAj1uRfEgLDb3C2ESmFoQa8AlIL/Qx7ckcKnX1q5olobi5/DVtPgrgH59atQBf8a3P9Uyg
r+DHw1a0RQjvsJAVCpcGYhwmI/5dpDTzFgkQ9r5cdDNW19i878OFYO3Vn/r45D3B0dl08vS1I4Bo
GktE96nLIxvbCDPr7QOJ978xAzYmv5ASL3tJUpNHtI5NH9TIIDT0PMERxAZ1866J0cExGE46jb66
yVqcoYyZO4WGHkwY2jD5IVVeeWNnecWyq/lvMaiGcjwqz4N3QxIgJ2q6KmM89X79bov7/UhHyZT6
57GWVNGc7sRJM7juXlagEf9wyoyiSVSrtGEH0r/maQhS3YbIaQ7/KDYUNKCsUyfT9WOIMu84rg8Y
qBIOJZMAjTYJ3IUJy+DoiwdGIsWKhA4qZB+wKjo7mhkJ2H2O9AsFu0yQMLZSNF5O2/tCNdGTKv0K
hRtidVkNNumh45JOWV+4Sz+ADaRn0kvoV+WKAzdjgZKlPjjrCRVwYXuRlX9yUq+V5VQ2U8wSJ1pT
qDHKVqo8Xq9IDqOWm9BuD1SLpCqZxgZnfL/sFZuVayG9X4Tz+tr5nrivA/CbYA6vbWeeCFOX6uNK
SAfkw6CiidZ6VG0/I5Jfs5e2PII08zJvLh+DWWRJYNJvHeebHaMrfHL2Ynb5DlJVfX9+WNZxreVf
lmuaPlM/Vhox6UZ1wU9Ky1CFqnCEGcAkEhKty5mEqYcVkoSI+4PAh0CkeCRx6OAWosUG+63aYEZi
BPYGeHMJK6iQ/Os/DKhtaaWHg9c=
`pragma protect end_protected
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="default"
`pragma protect author_info="default"
`pragma protect encrypt_agent="Synplify encryptP1735.pl"
`pragma protect encrypt_agent_info="Synplify encryptP1735.pl Version 1.1"

`pragma protect encoding=(enctype="base64", line_length=76, bytes=256)
`pragma protect key_keyowner="Synplicity"
`pragma protect key_keyname="SYNP05_001"
`pragma protect key_method="rsa"
`pragma protect key_block
xI5rRsZ8D/mWscsXgMgqvONi1IR+WUmvlhOeHpoqbkmGbmmCKddy2Qan/TbchxUow2f4O04cfAEu
JYQ5L/DafoWEAHShGyHztGxj4EyJX7x8yqtcAWwgcJlMfy/2Z+sYHVx4ASnUNZeQ8HXpWibYIZuP
FjkTNuAr1SrdQnqwhH5cviaA/5OheQSigRQCP8RRQlRyBxc+biSsCZMpGISZFX2CZjSyU+7V2yWW
ay7r6zDWmMmDZjudTCI4MmCNXIWpp/bhBBuYrBSF+L/5EsYX/jb3bbE7tKSBxKDVS/NsrCqqNgPq
LE6lSb2eW+8BDcfgsBxnkhOXEUv0U/y1UADlGQ==

`pragma protect encoding=(enctype="base64", line_length=76, bytes=256)
`pragma protect key_keyowner="GoWin"
`pragma protect key_keyname="GoWin2016"
`pragma protect key_method="rsa"
`pragma protect key_block
kt+7rNkOSYrcXqbgq36Tjy1mVNbqyEaJJcQomY0hj5jTsV2loT+ykCqTokaSF04RFimKeTBrbOMs
fGmY0J0Y3FLdb9mRm02LfOxlSlD1IAUzPqmK1XSR8d/4MtempkKY0sPLjad2NV3YwFQOuIgbOEwQ
WJexgoWi794m/yDoUFziRVt8L8gAHObe8TsXdCCkIFw1w5BV4qiVphOfsBcAFfGjk1h0eqKL4hHd
+knMywKT44w7gE4DaneMKpcCfQ4X0hNR6jP67PdO/EqqXFjgnAn0wypmmiFT+lBYDb/eP0n/hSzE
W8aox1YjaQtyA9zwXG2XZMpfhHFKcSJlD/u2/Q==

`pragma protect data_keyowner="default-ip-vendor"
`pragma protect data_keyname="default-ip-key"
`pragma protect data_method="aes128-cbc"
`pragma protect encoding=(enctype="base64", line_length=76, bytes=128656)
`pragma protect data_block
RvX6YNnGq/QfZrX3+SpkwDzMRMPNyB83XtyOs+h+gSiynn1XhUeSuYChhjzO2tVQ1rH3F/vCPrla
hD6VUALEq148nibJmMdYwv3hTk+sBmRcjCK49iKFYZ/tdhMSsIm1BIZrY8EQWICi7teBeErv3NJb
dWXAjbrToZfLhLs8dbOHQ5IeERmI2jxMHlIDLlxjLEHqV9ybINIEoYCUNFIKX8yrNAOSiB62AVk9
F65vgb+GThPHJp1sNpOWimfOv+/6Oo/W6BOOxzOHMKJY1us6t162gsKUU0fWBNrCj+vssOQq7SrB
crH9zn+iMCxEK0YZzuJkmCMWqZ7AZwtfRM+qEZNUA00xy4hADuAOa/xj7enRywhQzcafss6zoYIt
1lhyGaSALH9yhQlAkHYu1D0CdjsF2iZjIP5bXsPkxW9PLppuaiXqPlKiBsWHlmqTgUB8FnhBe7mM
kFq1zezqUIAflT+m33WmUalXKUHOqtdd0635eqO5k5eHI0wiUneaFAdCPFejIHyNFPCTvUsYCHSX
283+wbe1rbMZ+2ed6HIEA+kaaIKAxO0MLoXJGZKiTILw/G39+wS8OT5Xp5tAk5o2LnWbCSE+bBS2
gJ+5EK2PMHiPWhrKT6aXZzTlM7gHQn2cd7Jclduq5q3iY0AL5/AuDwITwSYQH0twu9KT9ez8D6tY
OTgXHwVBQVIcjZSk0pDezZfH41cqEAfu46BpbIxWq3h56AqwZ8x3EgOHLpvpSxxklNmRWyP2EywL
hh6m5Sfl84TE2Tr/AszoeaNR7okijFln5rsOGxKv+24JvMmMM0FSuhl2aSQBSIJPANY92jF+/+8b
d9vF8of5V+KIeaU7PAGqfuxhBlqWBQ4zcc1OvV3kUs3LxT1uBKtT3swa3Xja3JwFUolzJE/zx8cR
z7XR5sT319n6K4xUvhD2naLGMsQ5G4hHNsfQp2+wcSNfTtMsTxqiFGOaH+BX37mM5gnvUr51P0yb
yc/SNgXBvuBEoSNyNyGjUIFjxoLXekSooos7+DdzGJ8n/4NBrK693UFRjkeGOx3JDi5QqThVH8Kh
mJ3tELLl6f3MBhJcaaBUo9AHuCJyTtyLiS+i591GJajt24K1tilzt1/1PoF81irDg54UhB+6aJCG
fO4wGlJXfPVoFFbzGTjI4OU4gKQs0iLD7wQZ3GztTYB+E5MqY/ghXYQ3+u1AOPqv8e6cuGJI7m22
Qc+heGoOMGV1AIgCZFnNAOdnEXSoeS/QxnKGDaA8btg9SltrG/kVfInMjJkd3UvFpybzM8j9zs4i
gLSkVtdoByly+OKTzHRRPrDSoMtAVJ0JmXVgqkVqJjfy6DfDj5HrwLQQx9h5Kdfam4Va8FNYeMij
spsIKGWJ6RcKHZ40nDA+EXXhyD11fTbRhtOc0ui4+7EjzPQhuU/cMKeMSm7e+OFJ8LImQw+/Ufq8
qJL2dqTLUpgM7/BGpPcVIzj75dPF+fA9CELZ8hPE5l8i1ODEWil+6/rgkf7qIzUVCHt43ftXHjD1
F3Yns4n7pkm+hJ5xnBas7RRxixizD9P3kSWO5gTMuvlm4M/VjAtKqiQZQYjkFkTg+FG7I5rlSaIV
4Vj8GyaMp5l9TFTY1Bhl+pyN5PVzhqPDCh3Wd+SGQdgoGy9UKVGKnpGpt5978QaO6osIJpaAZ1Y9
h1qeOJ0WdB0RRjEEzTGaG1Wt1r9Rbzq3v9hMR4ILVkNqw4q+6krIiwTFgZvzRGjDf38b20MTirr3
R+dmuIMn9lgkadbWSBfV4mgsAUTCdbENmy1X1EMJLx9EqhCQkuCmCvZ89lAwfaDTIDmIc6oX/4Nl
UMAntgNyIF0s0IbrVO8xTbl4fSUohEGvrjpiUwcjgj1089urUr7Y0sCmZslzqBHwnKj8UQHp1PvQ
0D4AeMvJuSPOLCcI9r3UnwChSJ+JiiwfHwZLrlH1/hWe83+elsvPMuQp6Usw4HuRkAgKV+X2Peo/
p0N3EQaYbeTKu6usXYwNjwYFVExOeEFEglkhmFT39ArB4zweh3IhzbVfH5hVG57JUv1IlVHgqJ1i
GILU6iNao8AJRzB3Rdjh0MzFVsRaIPGwZ/P+pJMAaLFnxYVthpP9RgEl3/zIdDsyl5v1iWta6brM
sciKYIDuLPBH/hEI3RFwjFSZBV+5vW3PgPDY9DBZjH/FkWm0FDxWfsgUiaUdEMB/mk5113EjRgua
dD+8erOdgkK5E0zKrSO3c2qW9THrbhqL9LDQLLwzki8sWQY8IBvqvfU5ZK3VuJatFwFJamv50lEg
A/5tOM4vLCVq7Uioy1VjGNVG74uyMDU6vplCtNvj6r/9tLliEoD03dpoyeGp4URJoP+D38c/k3Lf
TgquqC/Vv4+3uugECDUb2oqUN3WoG8YEFq2q8xRIpXaSnzFapG8ygKqK/Lzdq16GOi8aJ+AXxlZ0
yHtHBBVt0t26tfGB3tz81kFRL5r1lpIEDsa37FHzOU0x+TMoZE+9EfEaQ74IYmcB22cF/AxD2ACV
W5LqvppKhDWzBDfOAjIY9vi/p+3rNRdq8BnfuP+33O2bQ1ZOa9FMmfoV95DmsnzjNyXrAvmdLBMe
DjZTBuW+ZWPZdqbug7zqveCmyamASgjP/uEiPmiUjHvyU+JYh5rXqwHDYglUNfalNetTq7uIIDF9
dTMW31JA/nwGhRKIUlyObCSkZA5Hbtt6JxHnWzlMicupJgDjhJcYkGrXBzp/q9UuUtipD0hraJKm
A2UKwcqmZGj/LK8a98sAOI3XGdZd9EBCKBV2K/NrLaehopCuF1Xot8de0YSAa0PIxW//7VAdR7fk
vg8cvOz+oGEsEN/UWHZl+XJFV8rnoqyZzh4kzN1shCu9S8kZbE4rmP43zuSNKT0YwJUi3pn7y/TJ
mFKmP1Cu5jHAfWX+7UfIAddCz/QSaQD/f/xNwm1tqwG7wQF+ihdrppGp1LGBtyruMfAzNRAV9F4h
PVbn3u//9W7dfnZNIwyX2D3qQaVDetQPdvzB88AOVhm7BtU7SQ/dsS77VXpmar6N0VeT+wSMAxzX
YsLIAUBwF8hWwSbm9Nt3neCwHGQIshVF1MS34/VeWjvAfOYvf48mMesdC8/WhVrPd9nzmhpxEvQy
Og9fl09m61W58CssKDXNkzWAOuuvIwXZjN1TFs61ZeArNm+6b7VGXwtvCBKVn0kjhrcgmAq3KcVn
Lbaj+UvqtjlCB48K5KjQyidsb8/HpByWozh4DVscDBB+GgLaIvD6Ud9iqWRp5zlJDu+oOaW1MZCS
fJ9llyWSBd954qT129c/N8JQn8doDnRk+ZEnY2JulJlxG+Z704IdmpOmeCN7UC1TP/BEzi6lpHT8
P081o68N1jH+llDoqfYZwMikFHnRSLz7W9TpvNRJAISpaO1Q+vo6A+IAMApA84Lys8x51FWlTPfY
SB1lPhKuK/abY9Q3kYp5hqhUvAIQYLVMWKi4EXSUXY4YRmCcethCsA/4aJWdfWgpjDfwFXT9IsI/
0+1gSSOqMcNvvsgv2uzf33O0rKmBQDpLzZ5X+FQHd6pHs+77qMDvtjly9iKFim/WAxoZ1P7Bzo+5
HpLEiFW/4AQMQDyPLXoYLBaf4binfb6zorydc6OJtuQkX4AewFc/HespwCk+PtBkGqfBDks1Lsud
YUcOfSaL+9biVHgi5HlaLh5nB4qtrkGOchINos9PDCb9DVK7ourmC5D65COGNcqAC02el0f0xJCN
npIutWQ1zUphJAPILXCMrQvta/AqxTZxREr69i4zexFNt3fXCfxSt4DCtua/3f1XMgEsYwLP3QQn
It51MalaIl9SOHMtotKC+U+asW8r1LlNyWLs3+NM2Gcfi9p9PMPHsc4mA+0ro39wBLgynd9/iAxr
VUFBWb134ESn+wOR584T2JHzwf97EWy2Y4eBPMueKZe0x8xkY2OgzkfNKOq27Qy8bXbIJa1lILLR
nmiQ4Zg6byTMKRToZwRBGejJuvnZXDQVeJ/Df4N+CNnzGiluzQ+bQR1HMqCNgDr1Z2t9faCOMCnV
q0UNLoH0pbkrd/FxTWT8bdNmLp//KARSZXivd4dXibAqHtBBdLyAtaGPRNqdwu2xX3xlKL2983KA
INAc45x3Pt/F7lR2HbzVQD6ft0KTxkOJSlTkJ7ZqvOM37gbIvLFuOd7P4FUJDaSbGFf7uddAPNSy
kmi4ZJY6vnKtyGeRex5vM3XkVRIKEBhd2PNW+L5vBFj4jd62lg/rb00haGNSNGeq0EDQGsqo2uMX
pLhpBMHCrLbEEUnqgLBQ6jkVPESeKXpraWr4HRbg6x6Bf6iNISRCyxhE3Bi8hkTQItOoosZ/hAoW
TNfKL6zU0YQiP8CfQ+/nm4fx4+BQEvLWJWzERJWvfeq7BKiSLrEZPdk5k8dLYO467sGD6jjeI3Ft
e0sIzIvNgt9VLU6jG7NiEFMzJKSPUrUZGwcfv3GsMwl4oYWNHcX5GN8K8jYv6UFxb8oStMRxGywR
TvAbsGWi96G5PDAhqlEBMommM4iUx0g9mkSfqfmJbBiGVUyCegVyXqvye+L25o226LneIGiKGA2H
DT6kGoedKMyFaNHmye31gzd0XeY8xsvANfRzlZYsuN+7HD1I58Di6x+aSRsjme3bm27AhdQHBFWR
Jg9/EZoLW2C1C1jwDNag/HHiMrKPAew0ZtLe6kFYSuEYrn0WDs6FmCcTpau14THsRMrMnHUOKseP
lJ2FEodPP3yVKzLWgJnDLG0Twfis1xMGb/tE3yfdH+3zeDSygO72slcsJNlVRVset5HlVysYi283
qfBw6sWg1hMA+9lTM6q+g2vN+2mHHdKnb6pBDE+lS1i9cM8DmCDYPJ5N/Z1TznBo48r989I8y7p4
5qDAWkFkLpGjyvmaJpEFWm16JGnL5DbDBkfBYzLBKhrDs7MlSywvgSZjjURnNma2aUGZ+nac23FD
1zDZI3Ue3YOhu98nFdDKq26Tl4nFWeaqemJXVFL9bJ3goa/if+LrkTC/Z3mKM2SuK8JN9q+mLhj/
q2M070/VEggYDWs11wu6kohzBXI4pP5GpaACPlaOBive0gxriAY+uoNtHePkY3biJnuo7ao3/aHP
StY1lb1iMHKGAjKEIqKcfRvutTfByK0DE5PQzE7ZUA02TmMlFli2OckXRenVMSgBX+Ra29RETQT3
hqwd7yKXTvrr7+Kt4D4ZW8+sybpK/ohp2BiG6ALnRMKC7dW/MN4MS8GTV9WcxYWfOkTt2hPwNOUL
hALbqvbfe8ckViOvJ+ITS1Q+1hA9Ru3F8BaoMbghtMlQ4tvXn3q+tsMpkXrRBOh53QiWbkcPLN8N
d6YE6zcE8C7TEAHfkAT6V9GOz7stUucrcKB0Ih4YsR1kuYhNxAB5ZeJmXRaZ4Ww4oiDktVuKr7Cp
RXPWc9yabL6tEpBUo60q85QeQlDOJVTN24vn6y5uno/T60ooRHUSGbuk2/mfra0wf7Z0x2iOcj7w
zPvLJ6828PSxUy0n/ASIPDH/PeWXDbaA6IJ5LtZaAHL/hEfaH05fqc9u/HVpYs/5SULaPJEah7NF
nw0uytoM0SaHqm+j4B+p6aS5HAxxTB3Ct+8wzyj63wpF3yiYQo6T1RxCnuDWCGhj6jQTiQPsoq80
lpd3QExYHTVmruhWfmWQQaqO2Tq7unOn54a7aSL4XBWZrXT/SA+/eRKLYzDE9Y4DonEXzUf3Zg/B
YVuFm2C4HACtm7WGy1KpnboY0jS7rhpKJ+mJ8Zco2WXTSKqzffLA4sULZXqQAxg7AwSE0aOy0dIK
f9C5gjX9xyJbsU+NPHgnBOYQGmdFx12gs5EsqrTUK6e+UCtKKzUMXB+0Kfopww2gCHfvA2ZSr20O
fKso7pi+pbGnzSoGYwX34aHD9EfHCGfYYiLcJLxVqJKCnqR+nUfRi5YIjJ5dSC9ESu71O8etNb3N
DGw2QFxsy7+F6EVg85s6OaHRYdraEEvoOXCdJZmIP9SPrmMPUbaqS5OiIRuF7qUj974brfuhhBf7
DbXcYcln+TnSw81jKiTXlAFG62WY4QxFH4xenKinNsKrYh3djnPLwCHnQYvwuN/e8XFLBkbJVzx6
k3F2kZq2a6z5bbNIbkZKqEX9Yu1rAHMHgm/5vflk5HhXdUK1JTCESQFeF79vmqnSWTP1eVgQ/6ie
vIxTHm0dqQ20929wzdvWDAQiTc4bwP/F4bKjSbyK+wrax7genguu7MNgDJxrXw460P5MsXMks74R
rpH9gaEWnj0P2npqGd5gCCoqMaeieXAS8R/niiqb+D60XSLTiiFbgIseZBLWeRK5eAskfciY7IXY
ViytYDf4WIA/9LabwbTXLrzUTOa8uII15vf53VjG2A8pm2otSuBGfomsCNQUfze9Cqcsgofh4Iyh
E5VJmxWQ8MW8XmON3iWO25n1yLt1PcjwAi6p3cADHlsb13CkNT7uEll4DGHELXa773ItUGN2PYft
7CXDQRubXfgCtTCAagMxput+Y792rAkMwxeAMzB143PLMiMrUMEzI396UkFj00EHPU9CjgqBlftx
syXDmuiU6MJvhwEIMFAxW5Sv0n9yGO/Ko/ujZ57Nqd+A7RPLweHH+stiJsTLve12RO81D9Cr85NN
uhwHeP3F/usSFih1Y48sUVC8Xg6OdxBOSs+F0oqGn5ZiCHIVkhIVUQAIAhQH1MY0hm807P9PifjR
xegoUP1F7NZQV9JHf1f17+fsry9pleiuUV39fGzRcPn63IbA+Me/jzIRX4X7DenP9c8s6/ckAlOR
6kd8Exnewd+905LkAqdCRQDEw+adT1OPntkKJNohiS3fqAZ1406QJ9XbrJ0nQCZtWZihYJysZip/
gzBs0eK0YMZ+yO15j0/OxLM2jBfqBaVrcWCrrwhQeBD55zaL9nl9ZybBvFWcwtzzt0VMHWd5IbaZ
CHGUSP4TWfuFziFH7PhRCMvoeN99dceUgFNzm0rMMF86/OeeA1hiGqwAA/PxULx/dk3Xi/zMPruB
Ur1K4uQDFnOLfe6+5L7aAvlJQ7JTNvqqEuwK7X461RNwzkd4nlfGm+kp8QI+b1gaOSW6b6tm3YsW
XpITQZO68nY2D8h5+bo/HPo6Qkxs+GLs4Di5Yasn8RP1PTgAvpGD8Z27dslq3nBz1+wrJHUozXX5
JQqrxAIgqHieGVvU1YOc4bnqGxp45N0QcGN+u46dRP0eI33q9ABrk68HyCawyaOGYjWVYKpGz6Eh
WxYkjYn460UwDoXSIPrPs2bVMk18iusDO35/I/hDIbEC8JV78xnFXm4KuN1+HtkegHfPolEYRxM+
SLUrC4ldtEWUU/Np3havs0Xfvyt+VP3V7Q+lO/T0ec7z3X99MWZFVhWpGsLAt6snng/5eDpYGDBS
J0y48fcGI5tC0As2Jyf/z+vXG23vSKzvBg1h5D/umBYN8/U2ufUNe88Jdw7EpYsXhvMcDxTpUNu7
B00xmZw4/vOOJxwDqoy9LXgb0enQxYvnk69CsF4EOa3YwfltxzO6eKdR497HlVtCsLodCV+syjjy
vH5c2suMmBQDX5oufm/DKRzVZq7rq9L8BOJcDDPfr4P2ExpT9lf2HwZqgHX/mZi5G3NdSizPib5y
0l4rr0Jk/2MGsn9gJOc7YX7HxnATWEedy4dDKNwmdRS01sxxNX9zVAXiRha9PlzVDNT/nzPFLXPR
nNjIeWw5D+Io9MeJMWifiSHIwF+CUJq+7qR4kbMfodCxIBjmft6ClJrQAHWKytJOMuYl2hnW5EvX
H6untRAO+0TwwD3Wwq8ivmBJ16x5VJDJtl5D5c9vR9y0jAU9ny5d/yLIh9On/8HvsBvAOVptQwY6
1doIqNLw5WqUTTMs6Fdr3mVbZQLP9fblLcF+Qlwi6yOdbnnv3HtjRimIj2CJQmtnwRVqHliBIIP6
XUMQqjf1q2ASlTPhx/bROLjudiN/I600KUU+Ezke7oiwsHK9OPl41Xwf7xy0tRL3A/EtbYXrI1aZ
RmpI2FmpM2BI4/axxaE+ncdZlGlv5rAJoKC1JN+RTlwPUt46EMCJhZ2TpncrUq1vvQE9iV4F/Zuw
XE5bHd9pF0XcooWxyo2/bpy/O5j+GSEQNPVMCxeMUcWI075otiprTAuJTvOkKBfmEptqirTaVES0
8nEF7oPomQqa93UQijQGJZ/Bs9rKvk+lhRBgA9Vglrssf8qjzkvG5cZbXpINh7QBliV/SV6a8zhI
pLVXvQztWp2tZ7J7lGn11Rx4CK9pVBFZvVy2aaz3N/w8ldgEdjQ6zZDHc0Toc2xeTAJXHNqz0Zg/
BNzV5KdJX3ucQgIyvzp508/jq9kypq2NFEfJCZqFhOlNdmGJ4grnk8xRp9gb4E6DjgVh+jlOHy1W
k8Du9WrN1W5QPfmigPYIBWQqa1aPv3xdWaXdIAlFPJyJzR/CeqOAS2Q+xbWggbmLincVoeKgMuKi
OAfvbszhjsxKMIfjyQb/gqUWKelqeu+hcb8lv8ofZO85g3r5Omph7Os5RJVJ4TexfGAh2CXNRw4+
1AHzMyL6Ixngto29L1k4/qqImEy71zFmkb2EHJy+d6QNrup46xhbqEskW8UrdSnoGcGKrn4kR0mh
vf/XdBLj9BEEA8NFEXxWBjcf/6f9j9RPE2WI8ijHKlJP5Wvfx+fH4PSJfu8SrbXBuaiyvPKep66e
aOpH7x/uCry98C/8Wa722NuiZZBKmaobFki0ag9xRkEdHzszbdLKFT2k5eNF2ibjWb6PzdJl0Ho7
RqiCwP6MEWpq1HE8HmTdCmvR8BaHgGBzJZ1S8ZIq5uWljyreAONTeHaxl2FlxfZj2va+n6PnwG7k
fQWH1Hq78upKFv0yC06seASCgbMe9sW78HA3t8qn/4utVDy3FuNvBgTUPeT3TirLxyNg2KNBojeB
2QpBsvqEC9ppvu/DuNK3C+1SCNV9r6NR8zFWKkX0r5E/72VfZvDMx0P/iF3DCe9+qCPWz2HYTWlh
oc6diX9EHBrGrV23Vs4lZ5PHS/T4QB7I6p1arI1zk3yZA/zoiowicox400UqOu9NK0JLuPAxAVu1
9d9PaycleIfZMRA3sCbfMb0tbszrF0RrDXboUlCThH3WdUanuU5FJEE20K7dUtHS4bdstGSOP4gP
cbcrLBZGB2LAPFLrITvRih4LAG0khQjWkjP03MfEtVl5GWwXHdplPJCy8PHdu7e5Nxv5K6aw+Y15
8zcZXiV55GhcZaKQ7p5hmeBf9hualxpfxHyrY3wexJWbAqheJtI106h1R6vjgXPKHOoTZ7BvbkOp
N3txlYkTW8nlkAkab65j4u1W993YflDv7POlNYDkswiVLqfWxwLyNmuP2pmfjuqpyCyzn19JOdBk
ZFehPZi8uCKcsXAH7V5WB1cf1KNFOYNXYI+4SLhAcOcMRmsQ9edO/F2k2irApNFsDqpFlsEtebMt
o4edBx0sHksy9FXYEi4IMI8n/FQcvWa38HDyMfd4Ifh7QZGIYWbYRHziyVEKo+4BJwx23z3/cxA4
YNe22KTKbtvmsTjmKLM+iLqA/8N9wtH/5gqoMjtCNt7hZpBpWOsclk/dV+A7v33cEttNU+K6q7bu
bJtM/r7YlV9E79I4NPmZHWVDBNm/4MceQSbWIZl0m7lhwkCqDYpzASXwIeQZpqRHPiZFZTtQ0+Ix
gKTt4fo1NdklWdAWZWz6295v8MDUYVKCOEK7feCA1cdJE+rZw2tonW0sEwcoRxxJ6erBwYvzb3Hv
iqSfeJG0nKf8MWFRo1t7Nn/xGKd9giBrX7jRvggS/3iBvAMFVhmpCeQ+Ma+0O/i8KAuscP7Zltba
02UPHaRpvUY54vbEswlv/sSvBZVe3lWFb+2BFvJN42hypvvPLza34IX1+dbJ7ChVV5/TQxBsXy5a
ABiK3MPz5oyDA0pfAE1shQWedAxFW/5ToEpLXHHttHwvy20jjcOvTj4JCwfgOhmpMWo2IPGrqthV
2uhZ8WdpQrCqRl5QHSpoWJ7H/K+/JALfRkxzI+kfUE3B+Sq8f3kpHbu6+bSiprb2xbqE/AhXbQbl
J7M/6akGApENZA4IebAKsfjG7i4RJU6iKFi0ql+iZXB4nMDyKPTIhXsf43+WxJCS7HnTimheQcKm
Ar2jgncWx9fyeIBfj9+8sufgQNd8vM/Azm5VPDg5Zk7u2BDGgq9o6iej5q0u8pLPB0BWMcfHhebQ
CV+jl2G4SyBRp0bU5kxMeRfAvjjbEsb6lDJU8ugA0ilElaTZt6sBk1ux8qTPUgAAGKClTQrovUF8
mNEjr8L9c7wWqV58XJbw7uFnlMWiRqzEYSg98WSfZjSNxe3QeF5D59B4LKMimIHWZM44I7W+LyGj
YLwOLeSL8W0Ry/TMu6NgGu62MGWC/gzEgeFNklJFJ1yZMqV534i40hWmpLzdHjFe6kgNiQVqSOBg
zsACU+JR7VHCW8vQuOLl00uFgZsaKuYphEbV35cQJtr4ZC1F0Ut82pI2Plu9uklVSKr97vK7bZWW
/DmxrhIGCTzdW0pEk7gHoFqF1UnIfsDEtpIywhNUlyj5O9UgbC5gN6vLyRRYWzFvK3tptbMCGD0x
WPaU91EiLkOueG7LgrwAK+WkoAQ87XgfpiZj4JYwBtJG5oMvmyz2e7VFX+IDuxXvUvvvVee4VcOX
AhNtNSt69klX2ODz0rgVhHMxLjpzbtw/raN0aZgWBS1UZrcxwlIuRP1Isloquiea5ExvYeKilkFc
ar4QVM6JoQUs/z9H2G00exRpz+SIpiKn3WMpvrkS4H1A/5laGQtM/8MvBir8yHZi2Jo4sDCkw4PG
UZiWGCi1aFQuDBNKRs/o/D7AbhMt4FZyaYGUxEyGclTqT01xPQH5RPtZskK+TpXKgHoFIHeQ2g11
f0eVHnUIFk4UyArW516AgOy1gs4+8Q3syrksLwq9UELfq7sFON8kIjXYtuLbnLP86jtUECTlVpi6
gdHxMiF8uDwxiSoD4eMeHZj+hyoZVfy6Y1M6EGH0larBqVIaKcjsgMpPT3+VttnVCXrUvJx3oX6s
+mfHo++n8P6IBZHugoxT5D6OpsA7alrciNBhtvyY8VOSpvV8tCC9tpXIjg5p5qg+BvqK1L9y/+oS
nz7iqbJ4jmFjtemTXNPwSwu5WaUe5R71dx89jkGhGvnvgQqPB1/enb1ipMnzAb2+hgn+jPRVz+Px
HhjrQjIFXKNLj5X03oH7EHTttnuqu+6swrdy2zd9EavV0W+qI2Mmnb2NZqKC2vN2WGvU3CtQLZ0d
3VRsJGkE/w0R0G5ksp4+D3zgArejqfeGXSc9jI9pdlTINoM0x5AZhhBZGAbh1oaBpXtKmzMrVXeo
am2goUt+aZdUMuhL7tbmDSMVYVy5pGAnznQHBgEwNgLKlJVVo9qilANkAcWCb28fzRQ//f9uNhzs
RkLI0Dt/+tnbx9l5shLHvXa73rd3q0Ihz5xhGw/XrOZo9pgtBnh57cGuVc0m1sxKaxhCaZUpFepp
QZyQWJ/ExSRm86lqGZAAJk5UgxQtldlFwpoU+LQMus64AQr6h19bR/klh4tCDt8KhuSUnsCjXID2
cQ8Ya0+yM8GrmJliWhgmFR4rOKcjMPIFNMJ55LyaGjyyTsZ09pQxeNcFM2J9+SRVmqifILufMX0r
NAjxcR/vyh8THWVP63ki6YYhStvGqNbQhbgyTqdt+I8ijKakfZUVcKEn/vxx6EpiHCKcFjt8JytB
N6anAs5vYfpQK8Nc7X/RoyhfIIVBU6QezsSZuaM8CpV6GX3EnqpXWOPkSMp6GVUqlrhEBMGp+yAl
YaAR2Jd7QGfk3/Fq4LHicihXIh2DEi7VCPMc82gCox6hQqkCIqZG6Laef20CEWvmQc/kWJb6sFj/
f4D3gURDut6zTnR7a8gStF+jPiAAxUXHNbqe1c0AYo+OJCaUhF/CR1rLhp6iaplsSMxND39ojMpk
anpDB0er1FE+G0/Rue1neGAu4WicuUtnFlNKitn6BQXGgj46d2xqHwbKcRXYwWzY8YE45tGOhfgV
IaV/DXUXvGYo/yh2U3fywmSxHOOOz3CnhPidK0u6kOe15fg3tX+3/iisPhA3kLBIKxgbjn19Ujlu
seN8UTGOfvxqs6/ZIPxfcZYqePrWmXwDYzysBjpbyEPRYv2afp+nB2/F6peC6NzzYdLNGXLyO80X
X9iREWdvdYppfKQjhhxpIHVRppw0zfNo7X86iJlWHzpyBacarR0ZmQaWayAAM/Baqp3V+N35SO5a
XUiNKV5xEyRopa9krifMCpsSUr+DARen8erRi89KyYipMSFr9MksTRUoIlgCYmsDTfw1jHKDNSef
IwF5IlSCthYXTIemJjPJMkwYOarS1hHWxzF7O3yt/dLSCCco4eoBvHwkRYyAfwzmFzFY1h6qt0j3
uVO6WC9W9nhOcwexZwPi1r6Mkosl6+gyb1+QV9G29+Xm4gAJtlLmHFgeAurjPH6Od5LI3xVhOPo0
IIH+jtjLGhEHGnbG60TP5Xrq6LFq1+jOAR5l060o6XKCqyiokoio8EBFnmcd+Bai+YRIzHuRd5g6
TEF9ET0BKPYrjaeWkN58T/gbpH4KnHPoPPlL5zXoCgQktwtVzQnWHpoXKvq/U2Twu9ybuPCBEOno
csWoGe9Rmr+l7puWshMQEtRq6e1LVnAyhBMwaxkTlATcTYSWf9DO8W2r7kA6wmtrLnHc/Z6F22DQ
dCMs4IRwXP6dCS9EhvvZ7bKgm7iQDsLsMJk7NpX6ziTKC4hJUKz7Qzhop2uKbQpcDQ4FGNYhHv5k
h7vxW5IO9OdQiU8RTVIezLfNwwvUxyJ3Dr3KYpY535vjVzOGamccpROYuf13XP0veqZqi9Z/aTAX
dUVkeDPNArqKB0XslbfpMizMGH1aZMnuKlSuw3IRUNhvxE1TdhkvC9vwGgbw3VlcV1HYt8oMeSrf
soaTrjQufn8f7e/yvYtNgYBThP1nR9f2Hjk+ZVcxQEhR/V3SFtyFhwPkP3aCKPffFnv2BpIo1VJ1
6bQJgcRQ89akd7bUGEc6m5KdubbK3wxS2rrJybSVbzE4ci1QWOQU6kkH4UKIpMVF5FW5yMOCuqxX
G1YvjylurMH5YVFdJJOXpg6CRJkk+qQyGb5uhPNn2yFVK+sUAD36rG/WVYahN00ETFdvU73iA/98
etByY7vSpeErpdiA0LWsRmX4FUNPvjH7YO96zzKuy5cCRBjAdnt07kzhmLfvznDXvyOApjMx0NhQ
RnTFzdc+j+s0vaiekkOZu97jUMeFb5WkXGOynpy6CsDev+nnnhhEs53W+xIHNYp7wTW5EKlkqk22
nb1GA+DjGPEL0WcQsCKBnqO62e4z/u3jUJoPIScc/gaKe+P/GJIsR0lGZRDRmm5Ld+tEjzHP42jR
BW/d7LmS91xlRq4mZmRBFFxKeJb4oClSfglD+f9XMKf8VqWIzSsutFk2EdVFDSbpFl+sgGjZQ6J7
Ofos+kiRmQiMp/sYGX5WsXICsFggPYMj2e356ztGVntWrjU+hcQDifBP+IZTAgrD2/RtqVROIJvN
tonZ4Ic5ZRirWdmo7cjb+fCZSzqhHwUkU4PVP0m9E5IOlZZt9Bw+/Wtbv4eilVBnFNC2DG7Z6cuC
4kBJGDQyUrZmHxuPhLltoNO0+VwxRI0eNLCJYaSWSVurxhNou6v8IuahlBybG1PIyxpifORPE/Jy
TLleBiOGOI8ZNWKId1PMwNLn70c1Xcktn78iqRH25pb2YMJn/AIcKbp6IXEoDAamommAeZZ4sRSs
UlLE6xPB+l3g0LdGO4bR5LKAzYHFLKSwBFhYfs10SaoIX+XgSseWP7oN9w5Idb6cXlTADRUjFHj/
MUae2I2tycfod8M/GsSqKF0bhohK0UVwU8bmWG86HuuhVVbRv6oMb3FW5Og3fJmd2vIP8QaiXB87
SLgD2L3rfUjGuVW+BcySRrY858K+xFCEmAB1VudT06JWOgDPlMKtpCAF72KcsWWNJqiOpmN2ZxN6
9sLwHICFVQuIYtPZMGdmoVRN0WXwRc5jjEuleoEkXexw3JNqZzYrlRBvfVEEsAUaEpp4AjizfOz7
A9c2VMjz9sVyRHpC2VHSOzIaFlLlCt1aJxD+KQFIf0SvQxwGZrlKbcPv/ITkN4ZSAGMnoq80pcHK
cUpfj0Gfh1iEtWF2lEVvfiON48G7mZ0L5jLBJY6/yCvHcHf/f2uWXhV+niLHH+uhEr3S+O9OTOI6
AvLqeSDd3Hkbxuiryf55ow3vqBFZcnzRibTN+VaNKA3tIY5DcuxShPfa+EJlxlF6pDDdZo6qos/h
DpiBGV6v4eR2hZHZfcelrJAZLSVy6BX7SUacdLGt93QSd90lYt6NT6A4Tt/eJWsp5KCaHL4VVo8R
Ym32OjoaQT+YJ6NzjvUVvmp6x8vQB9tfRAkAKma9Mj6TvrIs8jOlQXGcRr94vKUYzqCuUf/MU0XY
IyYNFH+H7q8Ku++eDSg9AoofERp82Q/C67nyCPLNFzIOTDCwYE+v9KjhpuFsYrOPqtAqS1fiLPlx
tVtctGj7BxMmMqnjJVp6VWHPtYCQeV1KKSuwLg1fruB/P2yDbQ5TqhFAtrlZxm+7JNfi6C1sQGLS
ujYsIirZt9emfgAvG6YmVbJKvb4mGljZ3fp5+PbHRwuvzlayYFy7xfDohCgqlHIBVY+p5zRiajpb
IEIi46RpvGqonM35UouYMxJzTVA3M9ciDFlZjsfABAnDlD+KQ80luGLsd4nKTzrX7zyZDlRlIWEe
gUsNIK0BTvDe7lS/w+nNK1T2Q46Fv+yyNqm2xYD6c+mBqTWzMc7yQYjNjRjxHoV3Favu7qtIm3lF
h+nEWYAKNwPwRPz+Bn3+DALb9E0yS3Wwi8LyIZjaHMLMOWDT9sBjUdpTaEAR2c4XhIxT2/ZYg3P9
Eb7j1fTswucWvMaA3DwwZ9wMBc+5purzvJeXvzZxdbZSD8i4pxmwCHwbcB0zxKrbPpgjrQ1sYxpk
gZPAF0F+z36NLcyokcN03GAmg9povVNFSOEYScXJBTa6O3Um5kxuxqo11OK2oOz/CA5Z9SxM6XDs
I7STDxDgANXa+x0Y72cv9F4GJJtDfWO/ED3XJNod1fQPKcAR1Ay5t/UADjWlDqOxDkmypRydMG1l
tkSM0CaoClTk1yDiEGqcGRbPKqGq3FqueiuCoS5QMOmihel8Yu0QwychhBp8TSVFSRr1b0Tj87V/
Pm2QgzfNWZWrqmdTOTdBo2nNNCwSN+Uj0P4AlFbtwgDpIC0lXmJfXofgCQS501fgRtQq6u7Y7zE/
mmzE6gZ2AY5kvXbYh7BMlhmSfoHcPM5wQmDa1GCvzIq9rnblS9MZeZPwuwocNWIQta003hoNEBNi
3kiPocTQueKmOzZEj2UJA7RV752iM6Iy2N6jM4NXILazN3LPGX83XSF1bk9TmGKYZmKavXHrsRxV
F7jjorH3FwwTBN2N9LGWQrA4lZ18MNUQL3H7TlsPVlDpBHghk/mmV9JS6XLtqbzvm93dAJ11OV3b
RFX59X9Rp/USUXUgV2Igbm6X0Rin2+Ie4lJXtrZiBToaARvikzFIDrNl0fHSfrYHk+4pU5T9rsGQ
/M3y2edV5XuyT1Op1LELv3o8TFxZ/N5bqKf7j6zMgdSs2J4Ss7SscQoIaSYraHkhPJM2avTgfGj6
abGYf3nY38zaSP3SgTOzDt3X0UyxMQkH20xqSFHZEorI/RSbuaJt644am/q5zbHiWVUxHhbqOG3x
xnZ82hQ4WItV+CgjGDz5U79TqWuUrCn9TFpbJrD6iFjONxOggQtn+GpNCnQPm7R8aYHGjdhAL8zI
vixURLkdXG87MjxiAK2n3b3NWkxKwLVIeTr7yE15t+JRP6QBPVoej3+vcryDSh7agshnT0WKG7qk
H2n5GtMpkuvejpiixsR0YildqZT1YTLVauuaJxMOMv9L+01Q9RBlNBHiIDPsW0t/QMCUXSFO9Osl
cDznXkeASoPzETD2eyZiRLOo1FsHFcNjoZcwcM3N1/aB7NmypYK3oyKHXzYj5kZZn9NjUrFbm2mr
22aGAyl98WPt9QvsGEs1Tjm7gGF0wgSEC61NZdKUtYD+YY+8yezGXIZmS1yiRITJNcEcCrnF8sJ7
msh9IukwxiyQUufSaByRRqvGSx/EWURfY/6MecirCncpaDPRfzq2/475X6kSCCZjdmqFgPbjywLI
9mklzzbRJwkT0o/b5qNML3jcaFOfIIXYs83eF6gmcPB98j1vHZziVn6WQR92fSJ01kWX0BrxbDNd
0ilnawadPM7h0h+Bwo48DfqlUz6H9kbZylCznhRLL6k+hyzb/CgDjukqNc/noqs+vS65D9QGUyRS
7odOeufuyL8vt2qFOWeDkUH+WR8IQ2y+LcVSd+oR1Sl097H+tyRkiFh0uEJRkkHa8Kt4Rp5x60uD
KdWLtsoBUflV5OntF9f81Ub2iCYkx2mbUJukUxji3hPaFpEI5cvJF512rvlmHEbcEYd6AtQX7hms
lM8ef3EvPEOirqeal4DOPbPEga3T6WdJf49kyhSqok09Ueiefp0ycRSZTrdL0u2comG7VNWXVisM
SFGc1hBGSHsgFAvYk8EryRh4P0HqgFsa48HjI3hpvTo/ES/hAuVpv+bjsChcesooXiuTGaGMLZ8I
DiypQIZnTT9Ia4NHTAfv5+GvGFxIt7o1GbrcKZucld5Un+qDZX+p+Yyqbq1Z79czYPGQyBTZfAcC
Fp7kqKaG+O78EewC32yhIU5uJrwL9w60L0A8PSKLLrQyafLgU0CxdHqk3ZyPhZLOoZsx4ChB0QV3
BeZGw69uz2RnqaRXF1lCXqtmzRUAEFP3z+3qFEloJD4nsl72jPeW8sdUSa1v6A+NvOpYFYhzUAQu
SKISCJXL5vPAJy/AcWejHfJSO30WVoqW2MO157uIPcbZIF+XJgqmn35i5ridWiMbs8rlxZWhX7OS
Fx5q7LKv0BEwRYvsV5x8XSGQ03ygqnRTkPj0aQRzRqV9G/w7mIq5gj5IZvCWfO5dxQmBlJRYb5zR
ivkNmsN3hUD2wiSXHTi/y5Jc/vvaeiDeQ60E6dcDbrhCrB4LtmQEoAb+UwOJnH0B4AsDdhgjFhlh
mO2Dwfr4Sr8x81b+JoHpdwQUa83ifutVf+LvD9jpugzg4I9bnelMsFYqGQzvLHMI2NjqnPt8ug91
xGn/X3tHr3/ZUOL8kFZYkn9Oy4kLWMKVaL0Re5gq7MfUeX2ndJj+dSXCl9Tqe/0Omzh6R7FbQVFI
UsdsZfl5deztuOd6lp8PMd2EHIB/BqWbmaT6/4xxw0LW1boBcv0/sVjo/aXfQllp/ki48DjTzgca
TKvxVMuhCVBATyLE5m5pgLG+mivtY+NrmvbwdJ+ht7U03V9tJBsnr6ab9ISbws3J+OdOurcbGsp0
UrD2h4T7LLUpz9vlLD/dpNEQyvwueQE4lWDe8nQ35w0r+m/KCjvqcmiHJfLl56z+5n/tAMWiFWuV
cSaEmyOrO89HyZbYWeHQxdXfCxx9zAMOZTKIKV4Ec4w3DKargh9bPdXRqosb97V0SbuiJzVHz6Sy
IHqtsWMTOomIc6G1Y5nKd7AgGnSVILXg8c5c3WlzCGpI6OMu0w3s+sAlSfO6y51yfwk2Ec+67w1Q
fGRYndioZXl57PCMv/U78TwP3ek6mrXeIKRvtVBOdp4KKnacspGCT4U3bJloJVPcAaN5IwcpK3yQ
IDBZ9rf0QOrN4TkLb4xVVKghX45H1lkoMmbxRRtPGulEci2oTazaCj4VomzXDvo2HYNLhZ7RfOE7
aNkOWqDB+find4kj90yPpGn8pZdyvYlyTXJN3qdr1lsDH9fnalPnbA2Wjy3yNbE6q5JtcixbPbj/
PraM1OODa7kyDNrcifKgObBgwqnk/txMthP/QwKDcQsSntJfESl6UiA7gaKm0GdlH98lOHZ77Ktf
glh0Sdc+QPrJuf0LoRDa7KrclEDgaSRHual7SyEFewFyHE1K4nIGvuUndaO23m4RzPwXXJRdtK70
1ELLxR/E/zTitZw7WP9DiG5NdQojvVe0eel6qkk/qYV5R2ZMeBwIdOoTYTK1lLT09ctkjlOkv+p5
QuPs/MxqxV2oLy6VGQNkybkTmiHgYlBQctK3d+hb178Ve6T3U9qHKvoplgxXBw+pNVc/q/pYTE2r
diFLXQd91fSIfKwIlmTIwl0kRYTWQKFleT8t+bJM1s1Uc+ebZZuiwXmUU1NtZYmpoz7kriJhctdl
qJH+YTpmuR8HxJepLbtc9mn4Ojji/hb6MK5kqUxVOJS2e4QHWgVuzRXxuNspZn8AOepvDQki19+i
0/PbzpRGqEUndOaTrCC8omc/zlqaozTtIWgBwJsRA0Zfunbjt3JYI+yzs0yaAEZDZ4bq8xkQfxge
jMBKH5NFAU1snaWPBoTnR279PMYqd5VLZcDxzYmKOhAwNvlZKQv6YV5ZUZ/FFzEj/Qk7xu0Y+MxN
8ZjucR4uZFrf9LmwCJwN/la2U9QBBqJlapE5iLl07qBaPXLguK+0wAQ2BvMqGQHfIB8EJItm57Bn
+w6pOsqndOlK8ZP7phWCI5U5iUhfnD3xeR50TPenB4VEta7ykoH/uKNS0gyd3/B/zfe4c8vvYCdX
UWGpjqjJNRxt7f4oncFhZXNhyWZj3nBIDr8uvNDgGExc36TPfd2gvyAIf/bqQTnWI9xuIh8j9jft
4U69GNd+767gv1T3FB4FlYLRRKYGLzkWgcH8ysaIgLgvE2ugSI8qsc+LxBvfwYRg6QNzNqOI54wl
vFJb7JUNbH1GUQ0T8MF1NqPTAfXBqivz9J0U7nGzeWPtH72Yaz2h2ifWa/UAB9xmDz4x0CdU3+Ve
qCDDEWCon1Gu4b8uiRl2BtJqaNLGWsC04E20HctrrmibUe2oSW8uCDD5rZ3CDTTQkKyfRt6w+uW6
gz2oa15ylDXmkFTOJGa8ETvdBknltVGL7+sVsYa5wkZV91IIUYCbyCrpPKYRaSoR1qr4VpqoK82R
N04u6tS3n6ASO1Gxh/YMv2dtYmMNpVhMY0AM/pqzBQ4FUtzR4oUSl8zdVeBnm1fxklASRETlSndx
qGbLpms3fp8oU1oNj47uaQeXhoRex0HKdjLA0DAVxK4hPb6rSqyUFZqk5Pw17E23agNzAKIRRwP6
vey//QIsVAu1O4sRavKpUNswAZ9BTFExl/H7pDbvUmvxQLwIuxsSkX61cCoShA7hZQSOGb312dEN
EL6ylDNbsDIOnDdtL/lxWOQ/4S1OeL0qokLwV7FvKS2vJPrbW252o5R27WrBT8ittEWEZKKfUM+s
DJZg/fFvQAQnlbMurr7x1RRUComaJR6VxvZ4lIExe4QrMVrNj2n+Bg/HlDIGTO528WIIoIwpf11M
v2TOsKkuw/RX2PP+nn1A+qdUCUGjp7D9/+hTDKUB+DOXOHRgy3KDGxUJr9zlwWS5aEa4DoT5s1qG
NJHhRT04Wc+wt+jW8IqEq2KPTJ/aXUoNg88Ji6RRKW2Sq0oNTRDyuggwHZl0kOWHwjJRBQPbh8uY
DAQCXxn78dKWVXUiZyhMnjVt2pZrqLbFq5Q/y35meDPO57Aa9nksqX6mtt0CDR7yCxiau9pqPk+O
shQmfko+YlsaVDMlj/6We8XauShRbyNCgbe2llRd1+kcHUOm5UfosBwbHqczpPMNFi+g4z6abp5c
/21xZrvm4Beun+Djfk8ICzy/eKEENYOVuB8kezWSICyc0CoFMyCj6EHB19YpJFvgLl/NGXVLEgdl
RTRbWvVLI4hGMOU/JaBV/zSZG1MlndZCPjB7wHX7G4s/OwPQI6781a9dL19MPwWc6syPePp7iytW
MXOvTzgFHNusnpEQQ49S0+lih5oyfBsC9hLGYJxsIT2nS1bf/nToM1URPpkGHOaZoys8t9q01BXW
Jdm3//YYQrhijH6q/a5Cky2agkrynuAMJChDquE9G1INifOA99cBIjQsiaipvGuWwmu9DKCnmW1K
IHI4eQhcC7AgODL2mI3fMo98iMnAPmFriPo8xPC7vehPCjIRbq1ErJrtegr1UvFdQ+smrYIV1YB+
MnTjr0Nsfm1MjUYLZbaQlNmO9mgU8/7YjSeHP8RO9v6wu4fgt9KOt1+cLpt9ejODUH3fbmm7B9oA
V9gam5xohW3YnMw7osP3G6wOa3UHKfpsaOOENfeEflpLDGuMe7Pgf257+YRJsVoeJ5qGcW/JYGNf
WMlSwA4vJkOrtgArAUgRzqUeTtwdWhgCdzxvTw1/6lE5OwqbjbaKHaTSWi4iXlqnq2nuPkHX9hlk
PCuUKvMKZ9O+m0A/2q1OjB6woP3ZOGOKDDbL7oAXIJHSerUjK801q6w3Zz18DstCGqdwbw/xzGWZ
e9cvlRj3EeO3+YxNpUmC82Ouw/0h1TDu4KXIoD2JiVH2rSiBFPjjYOk+jw/IfbLmOqhQGr/tpVJ+
6UZVWfftxZ/rR4vl7v5Zu5yp0EcpCsm2xWJdLYlDZrj8tDTsUyNB/7hrVTfSUnZgXC955ronMtCY
RyNFMhvyr9VDZE3CaGbyitZzxoGalRhlb7VCjld12rWDDG/7jqVi8IXaTBWpnPZOLcUylffSE/FG
jeKF2lphM0vai0Sux0ttneNN4DMTBb5+lLPZHumh68YjdHzJwZirdjes/PrH0W72y2MoI9njCLhv
DEk6dnFPK2HqPZYht/kfdBR3DgzEcL+CZbB8GaR0qdK1D8vOaqYBpoB+5OYhyObYUa1rAIMohc4T
SAhWErIZjEoB4M75dozc5LKksoiPAbXXz7piQQ+Dr+RbZ6JXcOgEMcTi52PsnzuH1SijkDWbSUVs
msMdLwmqm4J+OU1celgQDJytPxaQVe7yB0o2yPtMULSot3Oa40So/QfdZX2G+TuhmRlctlH7xBX8
MWbOgKkqx0OXhOvprBA7nuIL/CxbcvEaDrmzVyhmhpDoWQmRLedDBI1joMETm1omobmkgS/YxSs+
9aEelayIohFcKqgJMuUnEc0qWFO4YvrFEgjRiwsbW4E2HSCnLeA9/Y3pJKTN9X1xqb5rAL4VfQrc
ti2Ij9Btz379w6hwbhJQl9cO1XmvT1k8vuNdYk0V1HPBUM7if7vFXra3qZPztweDV0KoP6+dKfTM
08bHv4GHuGfN2+l45+ch8yiUQCyvOIaqoYpowIk+j5eUt/EzFO389aXLBYxswIAGZ4kv1Z7FqyPs
Yb+XP1t5H6SL4F13OukqiorDyxPlDC/Ra/hlXKs6HY1xGdmTpOsb10toDRrkQuNyv4W6j5nEuyg6
wFTJb27gbVkj88+sxWa+gvnGx9oKyOIs9uyW6f4GKMJDQHnbbavJ6irwLXAaeBrqA/c0ej0uVyVW
Q4kzg6tTTW8BZ3E+L7WrKS9JopEjDLnP4gwrnpGYltXO3jRq11czxX14Y7S/g5y5anlTKioGjRnR
Lr7+7of8rNHhkgklIXu+iyuG2byCLS2QPtZcQOK94On7EqLGWeKVWbhI1ulG6B2dE7YMKXTTdxLk
ukBZ5bYQmg57+zqkQIpfDgK/B/ReIdVY1qkRdIQsO1bicVc0GIeQq9xC0+WFRbtaYf6Jxfq+b8o0
op0pIekvyyVIR/j7Ogyu/kPfrepm4lDnEi4dxADLmR0DUgnFSB1b2q0+yMcTkEHsqZYX8Q4ONYG9
Exny3FgMNtDREoWEeSxHAAuLR5Y+Sr+JOVRRPHY7aL4dUlImal+k297nMDogi/XUTj2XshpovU2G
OFmSA5W7YS7rSw0aWPBvx8gc7LaQ2FsxhS0vBgFKl5K2lyZa1SDumRrdcG4fdRIbGfSCZl+Kgz+k
rnYK3TpbqX9MQDPKL5QGgAzWKshNpclp3nxV0KmZuUaumhszgClySgHajG8RNQ2xhD693Xin06HM
Gyt9nZVKUuxRMmPT3TTs9dPy+j0pNRbozMEVtOuYr971G5HZ9BN8jqpqVPOPLLb6sXwAcKE4mUgh
nLGgTuiMsSKC8od0Hx0SyJuq69vwyZ61N9h6SOEm9VK+iqRECUKEzLsHLvutIHVsMwqtXGCL8kpG
0ZJ2RiZRJ87EJMnObULc2zkkZyVTrWn1ZdV5DplIVG8mXp8qGPYGuUF4yL2DRbMxuC/Airpb6Hoj
HIOZDPCp82okqi6VCtPzyAxxDsoctovfJBoHEDTh9wb5ct3ILhB6IgOmFhkoVLFwXKxnxmWohLQY
Zc3L6BiIkQX64EXNHGrtznzVLnj5lngJX8cUH7xZOTkn9UpI2winyb0XdkRWnCKoipZNc4T3OnGQ
fE+adpe02L5XFZHD5+VjaWT9GFUYuaNroKTI43Qkw5ic4FQAn1PaOUMzSyjCM1vPuRdrar6s31Px
MLA1U7ubLXHS0SELLODO2Ul5NuC43hUw6MqT3UbdTZUrCXzhgizpTRn7SheX9hr27ycLHWyBSokF
ixL/CvwCbJRlUh0NKiddaajg3LqgtcZcYw20KqnRme1dTxtuCt3Z/ApvudJKD83HhzG3E3mtHfBH
jBw2TnLTMqRs64LitxD/MVXQ+TzVLTJoplCHU8gECBd998vDJ04t6WBx0xV6soCCUXlv4puipqmy
MMrwlazZnT3/+Q5AznEzJkDOpI0Fw/8XthVuUEtvl3yJqop0GIE8g97NiIIbaISk4j6KRETPWlVC
VqNrNdALOwwtlSgtbLyX2/t3aWkhNF9f1wlEweFip652YW8wSO7xXiP/onTOzVV6pzSx3fk7LX3S
Jp7FmPhXg2Fu/sg7F9c9lGS22//ePVib3OekeTY6RSb8IkRD3fWDZtVTLDdcweji+pH6zFKjQ7oF
42MkiI8oKpV958zl9byW9J6JbHCDnv1ms6oELHhgX5kbGJPSkEW+Q7FoME/QbkPGqGw42vPw7jdB
zDgDfsOAPBH3Qu5pNVzE4gmVZEemRyePqsZwC+QFf6hadkKHQ6zLw25iJsujACNBcxAQfB/qzd71
Si37lOcOrp5DYuvL2FwvqS/6dmWDYeG6QQB6j36npBkQC3QMGA06JIzx7qRlL2AGq7RtO5iYVyW0
V0ITeBdK1mqOaGLOeSZLxYOB9Tzwq+3wMeY+YDBHzo/h8Q2nhHtxcmmelgD+QfVwercr6wdnMpYS
vV5feOiNAuYJsQJWDGKp5qGPUaA4UUkvrecfpZe+0vgO1h2Nzr33+Pv7wrykISj4lW9tQ+E3ert6
0BaIHB5z/nl70FtGXmQCJZAnPB7cGBN6WrewdjuCbvtC4i2+UKUBCKbK/tswHOvMqN80wpRT9KZt
M0ozn6UrgnUgZfOknPCvoXSfYcsCAPs1aFvGBQ1ItsRzGr4s3Jez9oXVIb2NRd/DByOmECWWsAgb
vIdlWm0tnPUeUlmvc0ci+ASQfiUuaqx+MPJf7FMSGwu00QOrHzoAB3v3NqgjD2dzHc/KwPO7gvMJ
++3dcQ9MltF23/T2mBJ0KBpFeXPmWT0SVGpQL7KocnRdAthYM3bgUO3WRotQZogbvCJk8bgkfYEq
+8tlJMiOwqcWixYbExQ8vsbDg/UuQ24+B5Jyea6H35e80Atrue3P9kYMXovsVHtkAR5aioRUYmf5
TI7vOIYlPASxRwDn2UqqMDi3J0XuMD7gV/BuZmFYy2rRz57s4QSIlSR8pUI1ENKsGTUINRibQuT1
YOPWu7J/iUi0alD3LxDxTeOMowbycuYHQjcP/HEhFelejYhYCBy0MjlhzsAHvRpUgYW2MkpYTCBC
JuC+L3AOCPrjzBKkXoXojDhaBswdjP4pSK2O4wBUqrIcyv+G3nCcN369G9eJBPmhAki1AfeY7kRh
DsKZEQpv7qSoRXf3RJSKcnqiazqgLvXFS8reUVB/kbHTlv17gL99RgYnEZd/AaMm2cJHlnPmuTa2
y8+WiKEazb1QtCz8S25zGs6HbPE3XwpURrSZj94fgX+zgom9beMha/bJorwIYa/HdoWrqkLnKgcS
bD5GFbxeW0jtM7eg9E00ZjyRLa8ryqk6lXc0vFe3zL/cONIuUqM6t9jzOFBr4BLLcbZnXcETSou0
jwzWl0FSGCQGMGw0/wezqV9/jrmcRB2ASPHt8lHmqkklQ1ygP1lu/QBpLuRuGRX0v2gFM/R/1hqF
4O4JKDH0ocTk4l+noex7PidXtCBefienKPLUDMw+BxFzs0Elyr/MiA8AivsQXu2HiirPmmKx3NgM
4EJ5yZnmBucjPexWqFlcXGwVeDH/1cNn/MqOSPo5dGxBPygQexpO6v1DWRrjRsu3CN4X+appJm4o
w0PurLIY3t1kRSSKLgHUlRI73FqUyDiCCbsGEH26fHC4EyyzEF/m13suyLwQYxU8wMIfF4I7k+/I
YGr6foMas3FsWlRuNDCvMiS6aytqm1fhA9xqhd4KloeR1EkJgHIpzp1GZmMlFrrkneFpmhKcAvRQ
Yx1Q6d+UaSonlPFj5gxMbNF5nAClydcL9AAfttfM2fcu4nGAbQSN3hVeCYHuvCrphEE6gjsTCLDf
vggfhlksVlkQKOY0rTJCa4IKdezPpFDVqPNG4DaoeIVOxonkX6wMoLSzJkagWw197C4tJLmqddXM
+F0mrjt/smRGpKwwnpiRljMR1ygCd64oxBU85bDWSgge+88UNI8SGHF3wQjxylYM1O+HhTnIWX/c
rbYIu3a1juMjp0m1OgbiizSrt/qNAfCGtpkO0Oeljv5PTSC38Lsaox1yBjP8ctQbC6BwFNpCUB/p
x+oHufoyW9or2whSc8BVCk90/xqiXJV/sq0OurUfXZH3XJX83VhZ1b0Px2UjQ/FF9vZeFrcrIsqE
dAYKQEOZwgSV5e3cM/8xHtkVHhoMhPxAI20umZS+l8kVnVSTK4aE0tG5tAZhsUR7cJqDJEwGAg7t
vDFI81leAuJqIWMAvFidppiNsI+/jQ9MSVoJeBgdOX3vXXM1YeMXJBvXj0tWfeUiYyVOMjkr30ql
jOKdojyoBei+eLzyLPlO7vzPhUwxl474VaNuI4almwpmczmqdzOeG3q/iYvB8/iNJsEVPBYm6whZ
l3YeelJx/DcAftAR0yIcQqYwdidLc8NKvRTmuPoeNA7BWqpexNkU4LCABBER4l1SH43ZYEoNVNQd
t5s4QVtprvuDIxI2fRlFMqJ69B/ea1RQBMU3OZF3pUTgryjTq82iLCxOxEH8Cr7w6UaC5VSACSYr
w6zg3xfdgBj/dIULcqRbsrSY0uph0yLVUZ/LKZRpAxZDQNnCQzLXKY9mFNJ4WbH0MuDJ948l4YS0
2itdZDohpvzo7k1MzwCd+p09U8co/d7E9qqyWBbyIf3slBPBJ4LWA34wc5FADArmzAYyKnerbti4
CWL1Ft1/lJ5pPsdwDHEbVqedVJnmAr97zZBaOBTJ+DXlUlIQ/WWK88tFe6906XmBlXm5MCkYJSbr
G9XBMkUMnp8QN/nsOUdGRrztD+W6rKKf9fuNJJ6xvDu/VZ0qnWSAv5OAmUg6iXARN1eZEpcDUoGA
KRTGQdpmciaS2mV+ZI9qN9T9x8Etx6ltp1+vNWmcacoKL8+1DX8Dn/+7TeG4lGM1ubSeXuAnI9O3
gLZrkbA+B/nBXX78SJgty7fiIZXm5+RfCACtdhXoeII+Ndc02YYjDc99DM/vbaHkHLnf2c+QPRUv
v12sfhozQLefhPArHlK/L8EzBWwzOh33MQ8LmMHP8sTstvl2EEbx8VtFjRx86IVgTxV7tEzxkabs
pJyR9WEpP5LeCB42ppufBPA0JpUmohQn6s7rZL8othoXGxK71NmmMpt97qvKPS6P5BdY9DsMNVE9
avdavAhAN4jjmF9D8UGWusMLwr4gKVA5zUoMKPSIBLhK6qhbZEGvhI6QeqXrtAcVy5VGRqh1az3W
dU2aYUIg8Dat5thfOlh0bZZwO9vmizVFH7HeTBsUPI7b9yQPkBHPxU8iHX3JyVrmn0wkP2pzqbXk
SXy41rjJzULGBsv41aE5U3+iyjfoaQRmdGoKwOuvuvJvZUJWncrZMvBcRPl4M0QBKDbX9yYvLTAK
b8SPZcOIe0j8N5POsZrgJfzTSQeDeylzpvQPr16wi5fJVbiCTkrHMlFN4EJ3nXbnxftpPjBUKpW7
CU/5zEPXyjSCrodgffjmPMqUEFZl2/OlLwGGL6m44gc0P8Ze2cFTFPdewk2ho5L3qJrCgwaI3mo7
aGXkSt9Cfv8XQ3ZotyW3Tjeqxu/tPusYMMJ5PY7lxSZNeCEVSVVji+BDhbAlq8dcc/nuJXZaw+qo
mMtm5sYWpTs+q2Gv97Iquuzy44w7AQLoehSvk86p84zhzVPRb2TV9QK2EaSHJGiJfAMlu2wSDuht
fMqNonbNB85kweA3yYAb0i4Mln/DZBZ4KCzpNFkymzmVQVuYw0siMyKWmYs3E0yZ6WFvBBXHm5hn
r+iEdjUqgbb3HYsfhtguIkLPkquVjuDqZFfAsIrTxwNvMjATr0P4biydy+t9DG7JiT6IzQsS69Gw
AcBIX0TzhZbziDmpbFmYwN1JxF5RsGhhHa84u7jvC7HztRtUPXsEWK2qZtwAfQ1hU2jcBJ+UivR0
JyFRDdGkYxoqXdlpnCiqjuEmQdwemgbeJ8bauzVbILgkwn/R7TEe7nPwNYxJw4k+Ud/aPOZmW6JK
v5uEAto7DD20ehXHohgtxMa3oiqKkCdzuuMmtyU9mMXGWhrsZQnprmUqaC8Om5jLZbFSt2o2zuF6
CFBAOG8QxMHmr3X8YcpbQU9ZLfx3g2ZQgw0uHHNGtaQwFEDWhuiBpRJci/DJl6c2P0IUmPrzGYRK
RO0D0wrokYWNxpcZ8TEGxSMf69evg+aJx+GTBP2xmM1lMNP10OjO3uc//75WxsiMO+DoKlc/+6Jz
Y0Xos5tO6NjANzKP2GZYtM2+uxkAoTMHupPesCbcl5cNi67ELz81LIzpG7M5/dlikBq0V3qFYOkW
iPqgEzuH2ju6580i8ap4DhwhZ7dqSUyopH3kioOXdt0XA/4l7AWDWqs2G7Nbj1GpO9M9dD1/+Iw7
FyyhGjkTXPG50EB1ftwWpZw11+6RAmXkdAZRQ3tlQ0oOYZzqtPqwKvqroKef5iuH/E4+QKp8giO4
F1t4xopRMS8nXN+kW2omkstDt6rc4Kd2oa+Wq+pKKYXgFYH+dmNgaURPok3UBBFCl2Eg0QCCv9If
+eykdJ337tTca+qgIW8+vRnOFinALoHhydXPBQfc95+vLS1qjXJZs1dya6rHJ0I9SRHJJV2whgP1
xat45KTvvpj6qN/DXSUWYVBnYQI/VbMk+MUj4Onq98R/pbHk6y7ksuBbl2kREjCEIuwdUnFY9fcb
PCAN2CkHNA7nKL73PxmNV5HB5XvGa3bqwV2Glaw/SIUN4gpgADLl+4jiTSCy1Qsbog67Y0L4ICgQ
VOiJHDmzA7PO7YA2bXBd1tVM6ncD1o6fUhi9eh4kLL0wH7JMBXgXaZQ72QkTagU4lCeBi4kOZD2A
0BsaVQM4HLt7Ht26Noxvu42Lo/IqHLZ7c+yY+CEIyIwi258ioFAHqo4dhdM5Klf6OX0fllhD4/p2
h365jDfWYkqt6PDStky+YadFkvVA2ujpF87JvjtStiakhIQB8Q5ncE4gKgGbYdP2cUBHcpJviC53
CQrEvQjHa1rSjUq2goHhK8hFuCf+N3Mtva6m/hbBpwg/MGrk7aALOF7a9TC/U3qUxiytSOFuPFgW
0yBABlNczJKO0GNruoWheKBKKRaYgxYCl+CaWk0hM5Aj6F1JjWR0PvrjhL/oR2z9laI0rFrbxw8c
0enF8KoJdTPdfEUe9se18rlNvhdbNak6hW0Hxx0olPfvqguUbC+IqrH6TZHv2a2QfX6eKqM75MNE
24qETUG1WmziN1/ulasfTPADtw69fEpITcWqljJgP27eYRZ50cziTRcrHjaLI5g2mJN96e9CPBT0
YQMkcXErxBEAXonoI1O33xRqSUMtEOwimRAwePqwu1SamFIrsZ+ylX7VUuqB6U0OTLmbEJ+4TPbs
IEuNFKHxVVnLxanerSguRVpFvWLT29+I/EnRV7AHjYOVW9FdIIiEmjxe6717KK45q1QyTcfG1Fmt
0zEnkNItuW8RtSsh7nVG3346Oh9juk+cka2JM4ZfVDZ4LSx3o21lOeWcJgmpiEzczr28cGzMOIeK
tLXbphi13jxWhOtSNH/8iSyJz/3YsQ7KpJeJbHa/F29VrMec+qysQ1loCSi8OWn3Y7UmG3a9SSpo
AUAH7/a58TJ4qsRL04O2TF8x7FhYuXgg50ZSapju4XBU4cL03UERIUew7jWRUEAHCfqXr7o48Iaw
ViHOWL/COHKPfqsqPuAUPnzJkEtiJBF7vaYfwOLeswKG4ql+Dh8Ks+Cl2rF97FOBhD8jwZCdbBNU
9PPrtjvua49X4njqnYWwxssJ7rQc4IU2/ubPTAY0rKOIyRcRIpPOnaR2cAEDOVZT2wcWmnajI2Ps
qFtIz9VCyN1pmrGqnLsoqL0LI7vOtavynvJrZy4VSpByIpinK3jsdrwHgHzl2qoaofIXTm8/H57C
ytxGeMoW5NVwCqRaHh6TlvEVWlm21pcFTTeOt0n0WdP+uD+z8sTc/cKjhlNNHPX7BY5AkC9HFrlp
32M3RzT5/0SkuEYK7zgM52+UO6QpkhYR6Gh8p1LdeAQngSKfMkyvDt58dxpePw5FDZk9lEsGu+Gz
Y8BqP/6JBhCZiws7i02bFNSg1Wx8QU01bNNZlEisIHWKW20XaOqWOM3tAb7Iro3l6pSyk4eTUkYz
/gFKhsHnqMA5x8i3QfLkZVeskweGyf4e8ztC2GSpq8QPqMKv1hJWFMldEIxgb+VjHcNvxCucLk7C
nsmO9X/mTucuNLDt1+mPlfbneFpEg4Cg8g1o3buTXbjDBuijCES67ERas8uTaLLnMicQYG+mtSRe
Utg8izfpf5+u/go3nKx4cOrZes6AVY8ziWyRg5XNqVzwe+UCMR2x3mRiOBSodR6ppLgXPhY/42xq
yq/EE7lMdv2m3FYxQ9DOWAVHa18+Juc2uSkubQQrzTRUtJOOlip9xZBLicji6Bzjk0ms/5pJ/br3
6X0Wi0POvml10xfq9zOzCEBtt/z+v2q7hK2C9IP491qaIUcvHNO3yrTQwhWL02Q5b9roBerXguuy
p3KRmrRy4/VWZVT5XUWarpovbiJCJeQdLrXEE1IY8qjFnTJ/6Y64ZbHIaFK4Uf5FdElurtRxX9HD
lx+g33OtLkXHo8uOG4OZRBsaazPsExMGYadffZHPCiWZVwqJfn77Vvz87alLpoX0vvfTPKyrmDiD
FieXbQjjwpQH631esAvN996imLCvfB/swCczqR7OYGWIGoGYGWRZW60wqDx9Rdk/cXoNrwzDNFUC
7ih5CqESd3VsbcUYEwMXjjHcrjfaxEK1w4fpsG0hj2YQKRFOqD1gsjZ/75/xj2Yzkj21OOCgc2Ai
z/gEarLqUQey+3stlL4/NOEm6NYtAiitmPVOoNImfCPYtg7a34AQWVRJGswb8HMGdaHH2+b0g7s/
v9Wn9UGpeZdxUHZFVjCB+EkUlgo411hBwLye/LjI5HR4HivnlxQXMFtHjozPwPU678fqcf3PLJXQ
m5Im9SLTJMi4TrzRk0j1WjD6QZw2F/JFlGTfx1x1FH3rVOlhr3dgcLApuEkszmtIp16TezxxVDT0
SGUd/mWKUViQ4h0aToCguwAPHs7KLdZUPOhcwZd8rz0ztIDBufsbx5+RJlJIKYcjEDJk/kXNwpA6
7IxXxFL1HJ2NeHuoEZ8Tu3uhXTlXHdFwIl1jHTt1yPejezgQIxrnZEnDGPGRKjyr0+g33Ur1LTz0
rXIf1CyF/Uz2J96sCcp+aVep3P+a1Pl1OOi+THqn7mNzcsMikyh3MUlzkFbqi/RY3oib5a98xgNE
RU6JOrhf+3IBWwGeyVeQRisjck3lv2LEMquAk3MXvMiiGJqNf5UTRzdtjpUyh0sQob/t3jv7ExcT
1B8bsds4MD/p6+NEpF5LVKTqHOyiT7o7mVbgLRq+amFC8WF2mG6m6ohPtMcK9bd4DEOgfIsQrU7I
dOze3Ml3G/FyUNS8/PIQ5Dz6PHEDQfAzWf4Z85b7z3BteAja74TMuFb0hTweMjPIQ+u3J6EwEqiP
2H1aTCCQ0v3BvzzHcusTGf/epv2XgruPzCvm+Cq9pOBLyBj3C0MDK9SGGcXO5POnewQap08Rkh6X
+AEsrWikFAsjeV3X1E5u0nKWzZZmvXk3n+KAuRBYhXLYmU5fHIckaZ8Akv/9vwDeF2WYcXBb1aq2
bQYH1msJ8Yfl7Lofpe6y4O+PVhuC4aLtF0ExI6UjPR6Os8Vjwmrwdk+5NcXtA3F8fCSOkjeYrblW
MFlWRCuJ2AMGhImoELZ0iLXdWz5+ICUUfzmB7iAsLy5IyuyHHd/P4vE+wRYv/qMuszwBC5rL1+xV
yYHSQutcvh81AY+RW1MmbU0gDbybgqw9fqbxtUjbM1zzkEGkFZk4//wijvjar4CLJqIe/oUyN4D+
3/7r9BY6/9mj+9XddnWLHJRNNogKXWAW7N4dYH+uGVAl7N6nH8oCZ5emAU5SEnhPJHpLlJ4FEQ4y
BN9d0rJCTBK8gUN/caw7hw2nNexyz7x0NDwhcX1ua53joPC9NN0fD4cfo7iivxqV81JlO3lycNxa
rKX2/rKOFOK5Gh8HX4SlwAn/Bn/HE8fbPV8ZyF5FwVZKuRRL2wj84V5CrsiKyugzrJPNLy/aDgiq
vANbClpNksW+DWXttSbAzuB62PrJ1TBf1uPsZbcYQkX8M7zhx8l23l3Ia5DqBZ+PBcG/RMB/QuEx
ISe6mSKpOW5rymVYlJqZzxnXae6sfypikIGq+Ka7HRcJemZBJJG5Sk59fsHi/l9SHHGz5qHsf2Yj
o3e9O8KE7n5rImPfSjwv00Zm2/rBZQmlCxFOQLw7smuJCbdiuaToJbKRUsQF38M+akLAeb7FbOtl
z80fbGrWohiENqfwcsLkQm+JxKrnar0pEtU2E+lmHVRAs1FgXtSQjSGH/0jCz5SBrpV/RH8i6LX7
g1a1uRPXvbNySWPdj4bEej/9pKheD+9a/XfzwXZOP4HIHSjTx6t3FHAJV0ZQxQibbrcCGcibKKVH
v5Ulp5fnDoDJTs37ucGzOfwtZ1tzf5SapHsBV8jBfmdJW9MDjZheaipOfnB6MEdxYDzgDZOZbcjD
HBDhCV3TLrtZUG6not/Bwadup5tsEo4mgWm7NRZrpnXmp1aCAP6qs0Dk0N7et9BcJ4Afohm+Fw0i
MVneG8x3gBCEPkXdiELPzHMhHbjWt1sVx5LCWMUy8WI7lFPLZZUPicIrIFuQA087bSGCoA4wjLBk
OhGl0d9GXx6UxMAqiuook7SEofQrRF9CIJMvkxr3w3xtFd4JE4xgWh1+PNwjx4WSCmfc0wMPzbIU
Q/dkqwF+RYvDEdSmWkYLoR0AIXcYpHw48yfM7CTboGtfCMP9GxUXkO9l6YvyHfXf5ZtcoSXGxRXB
ZKma8ywchEf2Y29LgX8Koe1zmpQjuZsGWiGRQvOrpzdJikOX05SpSHz5xgz+NiTYto050GxEBarW
FWtnpAOz1NGpldxNOywT2X/PmkLNhbmR1cba8i6/HnD3h+qrXJBECV2t0WCZm75f3QpmKyyWqpEQ
DoZgg9cHCMd5rHc6VhP8g9IBxgAhEfcr5xxxkVqL8U6SYjQBbA/wkkFS604VmkkLZnfvegX8ytar
IfyPeyfa1EXvkc2t+LhV4aYVZeeeh+kcUBO9q/uB2VTNNa/r/1JzehGjBfEzUt3m1RtYvSSKEAKC
givZ8CFQ+oSQUM9NuUTqKPVyIiC9iFI4wlFmJAPmhlUXz//deXhoUd0jxU93ib/iLLgISpRQ0462
zX7QMPfp0Jnj7PQGIDLyVnjHBH343pDMq3sBrKDnwhHWbSK3Iy/f+usd6jf8Gc6xlrj17n2c/JCL
iLG50Cs+bcivaGOaJyO91x03P3y8PLT+RyakKp2J3cJ3WbVYBsrbGtvKiKytU2u7Q2dSLtP85u2M
0tV9wfHLqPG9M8VaYqIBoupPI1utD1BC5KkUffsC0pkh2+oVyRS0T1anJsTN0svrb9cOthHGeml+
rAIfCIJNLOk0M/UBiB8C8ZnEJXJpXha2HbiWTTSRSg6SU07h3kUuc6vdEAlM2mS6zLJCpmWCgSMM
R4HzQhKwfF7DfLXMcyCMeEjeeKQ8h8Yo3bpCPvmwi+NiUF09RIGwALtfHhLKTfUIWB/blx51I7nq
pkaWcx08+HOePMUJs2lFKUmTV784FYJmPBRJ/t8Bs5e5T4K44lqeVwpjCNCQbP9y0m0jVKlurh17
d76hrqqkC9GovMM02RsMhekxL6YiUB4nsB3QDGNE6i18ja9tLzLdIm4cXbmitId3i95+uNv6W9oV
XOWPIca16CRXSUGVI7bawh+O1vGjGbgP6weFwkEN7P9SAKZbuP8v6TLom2sBNKHbtk3nOJQzGjL1
9d95YNxj8pt6Rexbsc5Xka49iGExSyWqdgnAXCAcs67HVBbFfowx4iVSsWWYROwMzPT+r64zu8g5
VTmSEeo9LOISqvVkPG7/cLK9+qAg3Qn9xcRveDhkHD9jO8B3bVqFQFcQ0vmb4B+Wg8XlJZBLoYl6
Bsg5t1a5pHCrrX86qOabROZ54U9WkbkJZvyKZpUfcMHPgWCZC0aRPkPsmhw/vkTtKiExOvMlkuvq
8Bu4Uq4bdiCyYzX/ZJJanfOgro1/VQWJo4BEo66mfOZyjc6WogmRCWXJfmaCnQqDYEV5BjDrD+cr
iPUjUtKl2d0rGKX/9znMkmDeeaq4RnUJflSGE1agYPQdxTWgCGuieIhNvkHh5tcJCmCcNZ/YX6Ow
c7fRdSOyP9sVCwrj9iPqL+gw19wTFUCKK5lVjXaXCpiKBIJsqAmhL1CiteOkhlPtBszwlNx4FcqL
3MIF0rG/JKjgTcJCXx+LI/KrnOw/3XwfZZnBvQ5CvhS206MWEdPUfF0HM1A1EyiZzNeubORV+SOd
W9Na7Hmeck+KRzCvNmL7de4sr431GFLChU+uoPgcfkC5tGi6rDjW9P4lmk3RfFi8G8sCLcwUNp5F
BEjtMux3CEbKFhWFoZBLaxkuzsb7FnnoM6C6cVYq380KMbSVP83PUGbEY9VrBsQS+4Si7uUli4w3
ci8it7PrjgwVCv+Ow5gGpAMo6oKQolp9H4+g7XQDrUlIZ8jaDZj1Wat8Jn1urw8fihPJjCgi0bo8
tOICrWntjq3WfD3WjvrSiQJyQaIgC4YWk2KEP+mlDWNJ0Q+OS6AG54YMDgg1oNzAQGWYKEy77Jla
9/1ao804mK+q7csQeik2RfmNMx4LRbZY2+6ePjPDIhrM46IKcsjvy+fnqwrYiB2uIPPKBj8io7zw
SIsgX/c8aXDRIIgrMhk6jJC3zy7s/zhDC0pXJPIy/ERaKxKaSg953tUKngFS2YvNDlXEBV/fNyu9
/8R0oaTarM9PWNhSDl91xaAG4nhdCYGD9oyDuVMGf0l2JXnKoi6xWEOCzrZiGLYduVUCqg7URra+
T32Adsij3W64IZbiFnOA0ich2Poe1j8cktOFdfynfS932c16ByRGT3Ck5tDcZA8FLQ9YbBlFU1iN
rI3PFlgbp72vU1hmD4Bi+JgI+wRyxUwnxEkwR/NH+ieijQrGO1YQ2eEXxHoCPyO98GaAVUwbPA89
NfvI5Wd05fC2GTzO2gkTJHcZYo5PyGZCAUgKtoKlfTrbOX3Q3eFHb6U0jsI4yRFaVprjSmnaQP9C
HzE9KRCuNyQkyAlyqG+EKJJLdlXspJCUsLHjDjXZYZGYyD6gkANzY4OwzReKzZrbdMk2I9iJg6hD
eli9R7265kUbxDF5DQ6lLQkccJYXvTMGE+mbzWL51xj0GNKv8SrHcFc+nJckVOyQKoRrD/Zxcz4m
RBj4Hwh+XK+y8HuKVUBNOM6zE729QkT/IPfxePbOr2CuySJqvSsEXAdIjDwR8bOn8um9ZugaufGO
TPoIvhKjNkwwl7PL+DDTk675SzTaKdAj7cbHxURP5zqRghZw0f/fm1lWTojXgTQC9UTIn9aSaY+W
ccPAyqNZfcohKi4s8+MrjGdUvZI6FgfAQk85M/lDfA3yftLNnRQti9md5Xfz0DUGKcS7LkCy9z2v
ScEh2Fap1Cx+pjebtHV1g4wkPBxguFR0RZCny4pL2EWL+8bmHZqg9Wv6PGD5cl38TpWZQvBAyc2q
f27jfZU1dj/aLEcIk9BxyS3KlX9pbNkCVesqTz/bxgSLgM717V8fsafkYKKuj3iKTpJrQYwy/FiK
dC4eVEEJgv6J1/ww/83+SCbrfWvUS4a+CYBmMHUyqubfBKBv336aqtcsaB2+jNIEBcYWAeYf98BK
DTz+ONttdFIRsPeXtAoErgBmI7Xal3ej8SsAj3n/zb6XYdVP5Gy/5T/2vVtM+a8RxnXnQIl756AK
T8hniPtZrV3PIBlGfS8nkFoFdZ57qPEDGiBvkArW9ryGX2zVxFMibCQoIeI5DzFsfTTNqVjbrLSl
TCberFTEiKJyAe9qweEe8c0PdmzHG5/amXpJf88p5OtHYdPAxxp936w1RQVTvb8qGfckzeV3r+Dx
9xbFLjdoDxlfDheXhP/oA/G/u7YsUUfJdqibnYYju3gtQuMWWNWAmsKXCQdt/NzhIQetOEszjtCe
+e9LeAIBN+6RIuhJELNoYCE+xtm49vCMFaXgErVsLyumKBjykQjxG0kOlAVYFTWK9rz/0D84/23t
e7H8bycFuXHaD44gpiR5xuSfEJAmajTn+wGeyBaqbJ1Wy75n4pS+k4EZj14YDowi0UMGDnSc91En
YUMppGm2hj5YTEIVSqwcvy5f5GVytJkq/XqVoR3uhvONjtlq8qQDkGs5TtHm2t+dU96CruyxJNS6
HGRpZAjPHxTF6vnwBpbp5SxerCDf/378zAue8dF+1YaP4HqgDbdWngibAcEqNB48LHgkB8CdTE/l
NoW0FcBPGuoIMuW29bzRsmePmO18QCSE5NV/lR/Acu6Xb+MNJDsbvnrE5M30wblqJubedkVDAwRJ
6o7JM3DIhMCLKvbjHz0FZC/4tMQ5aN4q9LAqKQfCAc2Qj46miCVa/Ri5F2nhjFtmK/1xIrwUyYbA
x+itBNvbWELq1pGMVxKliOML7XyP9emcMgzyosCAx0KD6rgyS891jhVNw1CN2IQFo9+1kDphY07l
Otem0F0hzZCz/xQLuPTXujB4RbtkrUZwH2lEhseT40RLri/NoShcI92GCm/b9MQstBdNNyuVPM75
i+VMEuahLQqTKh8SglMywA2+1Q6u4qYPjRVjS7VjTLEX3GtCouh9qA1CeW1QaRiAIlvnMwfJuXQx
rxVNDKxabRP2xuafkIh9T0SsQ/vH9ORtVQSC6O3rxORWWd+Uak5JjbwvoSzSwStTGCbp9mJinBx2
4sjhGb37/9FNxTn+vEDRVfvlqdSpPCqZTa5ULtSEaY4XYDNPiUU0qm+7DriiBeaOTbY7HXlQktTv
BjAzYW5c8kde2PRBWa22yGdj1PwmhiXazdJT3yvaIIO2Ln1/52xuS4iAk5dNXJBTADoOzhSN6HUO
LMHtqYWdb7T8myUEx0Q7a/ksz07iaByZIcRlBAq0qOmlRx86ktozE4j1RcBdV4GLNWiFVpT8RWso
PlEtSdIkTMovkUmzTAW81oLsthFR3RMNIkPVgi7c3l2X4QKxXnDBCcLutvPiZw9rELj4v/tPXpxY
EXf26LLF7BHUkfJtCyPhJ+E3I0utmm2alZMYDI4YOUr0h8on8qVXkk8xpPNCSit97MFTSvqTtjVx
QxwUDF7DZFXxc84j0KdPJm4c8FZbAqRSO2n2bKi59LVRBI6TYTCJKyi38Dyr3dWZpYY+V7nT2R1A
cR62S11YXZYa+c1s2yKIueebwI/cHnCE2nGnhACFF6V7OWb7vgLw3Gv4iEjDWj/3XWKemDVzPzns
ydQyquTD6W5qLEu1f5Wj52q7UvqhJVOd3T44afrHvAMuCdrpw1HxKlxSgi9v4R1akN+eicw2Hspz
32O23i0/HELI/IQd+MbCJIm9hWbOX2BGUhPTIIImbY/N0xVIlc9u7NdjVzznSRIGoIZR+tvRWJeb
+iJxiUTA5UskLYr1Tj0L94YLbceRAFXjsmiWzEsUvqSrMbyHYIB2jFhenEb3AjWGqoNmJBdD8cfD
+sHiqJInEBzSFgjx1/89Dn47GBp9+h94gF2akQInircTN3oZX8GbD70VeEXZwLwMCn+bKWT6TDhP
n7np0YsqyjdqqzgphM9D+v4gnv7uiyzYLKT4gOxM/oFZYDvIAaXnXwrzSWWA4vYLRSboWKb1rHJY
5iDqCutIqJpnoIdvCfD4fkyVvT7oq22J9qTmXw1D1TQFoVPrqJ/ZJl2pVYG+oYutENX59OM9rM53
WKIik73QsTdt61t8g4SgoBfT7vGIJ37u1XKS7iaLNosgD0H6yFXT/SLWOQz5Cv1M3Ys8EfB+yfz+
/jceWL7PIEW1C90uuEZxsvs4izsOZd9ob0ZtooWxtzdkS9uFjgKJJkIEm0Bjiao4jlsTNfKxsDg8
iczNS7AKH+ZMmS934Dlz0EI8ruAtfLpKH+ryKAJqQsRtwd1gHZDbuI8KFxC0YRKXZuVoA14crDvI
+a7jvd/17OBXqaw/jGUmSHxWgdOdFuBgYCXcn42pOgZFypVo0ssn+AE3c2AHjhHwYFW+HmsfxX6j
oLUE3Ocwls7DlK4PzJxkXRQdXnVK4s0kjCyYUfedhhSGnJhsPcl3t+zJVlBij47GuyjksBJFFY9g
E7duqg/8GMwM5t830PlXKblX2h9A+eB7Uof1XJdKIA34dsHAdNYSIidN6sjjURPh4mo6DldPLmEY
THuVQ0IpqrX2wKNIAJRG5N6ud4jmqcUCicWvaoMfU0aYvwGUDERCYus1lHy3Nlrr+qMKA26OHJQN
sKqVuoYX1KmJwYgjnjFZmXoWzsJ8/0GEJ37vR/aP7GvsCi1FPV0EMNRuq2xPHLfVWFjog+inZ5OZ
SA0G8UJ3tBw8ZngPfyVXZ5ZAnQiCOiBw/nf5t0KYTj+KfzLhhF8IfFACyTMvWVr1VGkx8fnu8uP3
QUNZxwZn0aYlfxy03Himlgf3AbcewPRHIbmdkBbrhHp04aWErH4XeIr5yJYmLb4AU++UjwRfGye0
GJekX9qgJiEo0PeiN4UhoazmuSp8kAYxlrAP8J7/zYNPZH9P+DTEyhMFNqHiRvowxGF1k1P/iBib
k8hmno1WxSDgkm4Ov4j+PFY+BDfPujPtmqF2fMLaG+pvmdLwlj3kGxmOXKrf7s3ha8bz6y0w60T1
3kEXHD71Ut+8aoFMwrCEmBjIdfgrWwW0cOT49ELvOlhda9VAszE41dhbiUK/dT0/kVicK0Nh4JqH
zCUBuXzS5JfeiP9LQp1esk3Dbl4zEVMZY2zCaCfaGq05S0OzB9aFN087CIz2jWUBKzpd8pRDSj68
WGImPCMPi9SeD4es9NqM0EtKncTUDqZcXBeV9gIih+3fAC0bkAJQmynu6q2NdQMFzqR3+suAtn7F
CYyjYBOZz/WZncx8L6d5BzEHGrUZRQcQmWH0WGDOEGRcoDUYm+Y8YAha6QaZziqYx1rMincF5q0n
Hhs7vHBlwxo7oy5RBnKa+7rHh6AcrMhWmijc5Qs5n/fzfM6bKRckMkFQb2ThdpJ1IqN0l73zJWhU
orEaRuNIxVnsLmqr0s4sD59MQ0F9D5A1UGBwkIBQoPTwUvefHGpQ793o9kCmPgzbSFf30CZ3QbhL
m/0G/pjFErKTOxLecP6wpERq5B0as5+kU1sJ/ADnm2f4/1sktguMCbk79rlLbrg7411VJ6vuTwz3
jpynZcsD3NxNISCJoIOVZ9WvjoqgpdyqbFSWUDBdG4stO2oOdFAUegmWDqLCHEdsbswOgWbYFE5r
eR5j6p5L9aY5r6PfhF3HJRn8WHaujs7FuP5w9LYVFR8cYKg/FOmpFWrTsCEG0gKpyyZnC9Qd2c/u
BTG+YSYVOQaZFVMjf8VJfXO9BgPsZtRe3/tgg51wz/wvmAZF7HWg8Pjonf8yi+LC+T0Jeht0rmG5
UBniUyfcSGdFi3ao5g6xrVn5yCkPHAP1HVBh1Pv/q8zukPiKgx80okaHd7+wCj7gR58y2qMwGyAD
1wNbc7uKHqrGzYco9CfwtIXov/5S+sTb8iVSle1yYTNDZd07+PbjMnyeu0xIcN0VhO9Fe6A87Utd
t/c9jHM1Kz2N/Q2F5KTHYjMO64sQQ/cFY2JFuVfp4qY1h7scHOdig7oHU+K86gaVf887XFDkynRG
ueMlJ2zJ48c4+vP81IgIPPuqUt5Sx91A0X8oIuCycDJGia9ZsfXG/QLKZz5Z03Co0hUdGOFcLg4X
1uuLG6ftATHDBnfaiiO0K+eu42Ww1UwlMvk7JQ/cXU4br8kSr6E/Z7gXR60ahpNtwSQAvwC3xaWn
lBp1iHm2DELrqObmTnMKy6dm5iM10wQQ0vWOSj53rrPx68AeQP/4TyYGBXW03DIkDJ6KabkFt1xy
rxMyoAH+0iOemOLMPw7KxY1MgHZLuN5cIi4add63tWwdrvSADuleHnrbKqli9fqX01ucN3efty8r
dMJH6VmCrERwDfqrZLyjyatnH4Gx+zn6qwewGvlcYoQnBUeoW6f/b+LlhRHsnC6I+Lql3E6dY8na
JcUbm96beQZSONCKICCYVot3sBiJmmCf9ej8y69WExHxFurhnSdkiOdgcLr0pXDXYFkwfWM1I6Ei
WQoCBYjVya+vlXFyOJPp3ufDvBopDeVzPdIyts/YaFJKDbJBzSNwQEqUSd20tMSjrbxQdPzhHV2o
gPhGoDA2hQp+/DiyukyhUbS9cl0lX1aPTDkC0pM9ZCt7Cii/IKph58CpSghGzOwBMjaNkismxpcl
qHt9CXwRExh48abJriiQUkQ5krNcsEaHhrIXwMDDE2/Mf7o77Xu728XIWL/m4FqUNt7hp1f5/Bz7
hMiRMJxCaKWr2MewMYFvHMtIlu6+LK84bWp3mvh90yfWUQBaUo/AyYF8HrPmwIQoj2oohN4733Xa
g6FxVvDiJVzxs8oc6wpWOY1QPG+UOZb2lTpH3aXG0CXF4fp91maljlRXfR1BfFPYC72DXAFAMPPx
+kp30QoSMWJKfj1xg3nD19/hWwJ08t+Nnb9vMzOV3k9JpkNvNRVXpWrQczgA/+/CE7Jn6PnwHrxe
27vzdLrcTDrWbzDBvsG3655sbEUCA0QBh20lPh3Zei0Atp3x+wGA1UTZQEs0l2DdX5q5s5BFdAQw
R4REiDZotbKPN1ucxS3tRtyPOS2UXZJvapz5tkspWHjsIAU63784Q48mJcWSHVvB1zAs9pl9GO1Z
bBr5SW6+Fj7X1XPq8IcHxW82idSbbWo2ekHbpZGp4XJREW2WLIeAs4ebS16E0IARhCGkiWElVsIA
iYyjW0x1xmkRv1raGrVrG9fmWtKrNv7cnWnvNqFWL1FAtPzs2tnkD/FrRo3vUwA1Xqv2n0OwsvvC
zayXBgzMJAfO4EhZnBSlXhH/i75NlP5/U7l1jwFJVfh9YqntiMaP+FqH7KYjHaXqoiBF8ZCP5Kl5
5DZtoNgng5Cw5jz2r3Q9nT8XTvpHjUEkmqgDqUwtuqI32v2G2bLQgfj1qrKkjPnnmIM4/pKw40Ix
/DapjjA5dV7b7r/WLmQx4IkHUPLu55YeTuvUHtwwaOWgzGzlU8iA1JQOkdf9TSqzMxUNhwuDTvDO
0xQqPiP+I10FZNqbwMOhG0YF5/Lvfbv9Ie0ZVTKTq1GQuuvpYGI4ahHBEXeO/SCXbyd5eF/eKKPO
cOBO7dwUuXryMBrlAwuAd9U4YznRo9Cn0w3Hgmrp0v9yp/ZwrYH5OggdYxOiGuauKtRHofMZQPV8
BLR28w9+zRUA5+X1iIGyJ6hKR0lvqLucBMR5EQNnwE2Nc5wC7/nozBdtMJiFWKPRy95NXAsgPT72
d47gkk+nsxDJsanLnKH4QFdt/XlYPKS2qf6OwJ9cH276UkJv9zRXFD5NzSuNaPUycFwbjIbBY6hh
l16kRsiun6kBM+08epHAxUKsh1L1PYMC1m1AGYoqFc+uflY3l20tVyE24fCNUzLvEqJSNAy0RW6u
8L3Pdt+lA9Vs/v7gxYhWTi/pGewXzkBU+5bbSPMvIZ+zQOPTACevZ7alrMGDdIB2s/t3kPEnyI89
V3L+GMk8SRfXjujfdgswmT3HC/1PimWCE8GgT8D75yOFXG7CB/+OK5tWCcogO0sYS0hTJA/Mss+/
nSL81CtZAh2kfJ6tuy/VfQhVPLFkA/Iu17m5fOpnyvHbOkPs3oabisDhXGxNFYHRPeJEb5o7+qTt
W4A6guGdrek4MrvlELR+TDfiMxhySSvjWmQ/Qc4xi4YB7mcleSfEqyR4pTXq0MFK3pzSdkYTVMG9
9TLozEtU56xjr/KunYbHSYZqa5s/45ZBlW0frpjcx0pKyaGHX5fgZ/2KiVccwiok3ltaT4tYxxqp
1ND6PF9nOUl/nIq24Os+nYlDSPQ6+edQ8nCvCi5t9IztfwdqIVh2QLdU5IQfouG0IXuSp6Bu031j
bsfgG60wWRvrewLJA6Qlix5bwcYZhy5npWQZTgmdpjAwoSsucepct1nbaARsDs+awxltGusavAX4
7YdKSVl7trZu39z4nzk/w1zwzJMD7fafpJf1MELnZzLQ5jF8JkJZ3lSWTwG07PzoP5SgWz1oIaKi
1q5E52HXYIMeG7NiyOkZqWHQtcBq6sO5tdaiGIC4soBPAvoH3WVQd5KG0dVZsSj78//D6bNH2smx
Mr0/KaKRjby+a83CJTRm1n+cX4ZXZs23PWRSf3fTSVZzwE8dbBUlFo/CIcuC1mCoUy4rMbbpSTmN
ZUe6N1+sEopYb+RlmvyhWp7jH8zisloBVEJ2T4YEdmxvjLsWWC0ledy7tQDg7Qw16e3WvlFytANi
EPNy8dK5JDQIS6EyJVAX/iC9fTkWiGigX/IfceM27Gx2nrYYLTQgSlc7zHdKuSJGVM3YOdotTgIh
ygxrk/mJViKWJ5oCZJaT5q7YyJIgPqVK7L4p29JPBqKTlIlXNXq+yXfOgvwHapPCeUtevTesKlwZ
KvyNF2kaD7l/14/V1lOeX+iGBBccnw08XVYgUJ4WQx+BXfHbqqFakfGSF8hJ9POrjMA6zxgraxjv
3d8JQcahMzdbgJKT91n6eJxbj7ff5fXf/ScnnyJRd1swtTrFKPcxnTYJwfG7ACJykitqe91eJYyG
nL/vk6gPcqEH2W2s6JPFrJPVsB0ckxgCWKwXUK/+pG6UxHM5iFVP9q8Fm6rnmv2w6oHrO9+t3Px1
oFVE2gHSf7K1vINnKmumShNcc59qkgB0pUG+GFcVkjsLit2q5ZuFf3MeUz+urPbg2uj+xssS3YlA
/EvdE7U5bXzyqMJZcz8bgSW++cMKKQdnSajJTCQrCujwM8D21tuyji6lIbUOkLWGP0h6nEiDzmM0
UyeTCLCpdvx7VAVLRy1JeNHArxDeUilB04SkP7YeBYRC0TenfRfMiF5KOA18AeIJWLTUF9Um/1y2
WihYpC7NRDFSlszgqqUSc2K3ybPlxPJ55vy9tQVApRXZTPJUsIAQGhA7FVaCve9AM2l9+a/ErqvJ
8wRC7TNiM5oYhzdrYMZZDQ++lZxsQSRXs0vIlm7+Dzv1dWSBg4rm3LE/6hz+j5AyYHalugPz0dQM
ukwz6f2OxRun66yzdAGtP5Ef9lBlJIgiHNB6OPP9k09ebsobQM1FAVIvheywLrsQI6A7mrQev9bc
S0bvcKxD+dXd487+RJuHvmYrGBHWcNi431Beb9ly5ItxiWh7RMNwxghfjSXrP0OxaiL8Q8aOlXu6
riqjTScUsS21DBDmIBQf5keG89w28Aam1DOCNBt7QtHaONa35CfQ9sm7x1yvWRSolMYDkIkjOWjv
q6Tl7q3gx2GhEgFERprHCmCaIgEQksURRmoQIuzMGCVozNqiK1VSnydSjlrjPJo+4VmIdCzadULx
qT0qXhtGp51R5yMJpQJ0c5D+qqqRwvf/5vQmt9EoTF8yPWOfySEQeNH1vD79VcnxXxvT7Wq5kJd6
Lg3lo3PJ9H6UihHWRMWH2xAyoshX4m/i8lnlQWxGVbTjaJCQ9Sk5tWA5RNEakqBR30K9blBJEdDJ
K4YnstuJO1uwea7kcsVaAtZTdZ6NaZAfzNw1IyYcT59rTnndZXFJY/1W5PxyfACjVSYWgyUhQEOW
lFBJmisPKn5id/+WcLvYWVxL3pUV7ge9hkpr5H7BNtQp2Hwu4UOksbqeKLFsdnhq4+PvsBhqLfaI
1jA/Un6myzgDHR/5ylzsDrhrATX+AQ64f/01fIlVl4Wkfz2epQthlqBqj21+taM6IYeObjJMVQyw
OrcFHvxHmSc5W2fOZEu9fX5Ccn5fTw1Nr3mNfPpwaiJ5c4Vja0RYqAqtRf8tweeBLVQlqkHVAIzT
ltGI8aXfLdhru5LdZw+mcYwJfuIBCVja6ol0ZyJH7kVLcabqg8gbT9cp31t6b23VeTGXTmJYEYRn
m/cRIWy5Bo3j5XvlN4HRKkAMFpztIuYn9yJ/PMpRZcO9q5+UKVdupRFP7qqmJPECSRD/UmcRgUS3
4vW71rTnOP4nN3vdG2955DHOu/j79OwLSnF8H3tUmUZZdI8yDkIPFNAcfrA0YoemLuz3BMDTFv34
ZlFWrtRdxY8eHuWv9fu3W6A51MAbObZPb/bRBHIRY71IBMgyCR5YAmi0V4z1ui4a12piQ38kL3ez
viC9CHnOnYQvE+HH2rJXMfSh/S+3VozstifHLUR/m8SdlPY/ajIOw3QtgWquzG6E7sMM+R4bgYaZ
fntSWbdTx4toD2scuBCI2+lN6vD5gQGt+4PJGK3c13gUcYw3YbDHeN1X28fr9jIbJlCm2gr+Dq8d
qXGSU/V6iNLbET4chqUE28SjkkIsYIhHxCcrYWzMepEedHgTiI4SyQpgEm4cNvzqiC+WEuJ8AXbc
7XlEbcb4MpcE1ZL6wJgD/YkGcKh7wEkaPQ2r1lYD10c9otwpxtcIuOb2D62AEnuYRS5Gpg52WK7s
GTCpgQRspLNgJQNs/Jr7gAzdq6cakwk6j9i35HoBIbaNUO6TtORVwa8qoEg6jsdSPw+zJ64EWK43
z/cYlf9klU0l2q4YyBXkMXNoRfRHj5Y4vyYpwCsGXvn7jKL/aJ4WSr1b9qqFuEnrF6PACk/U83te
uQN8CCBACjDph8Uc/KSDXFvFa1VxhKiUyM63oqQakxgIi3Xd1oK2qvD4jH8eNRgz2TjLbuZZLrYb
cwAl66ResapPzynEBFfAkLFfZQi8CmQMc1JO5yhYdUrm9pCSurl1tcuYeRNl7vsDCoYc7dC7u0zu
o3JvLhRx31Su41VB72UPQEbCbjF63U33MNPgnmFIbvFeVCURfjMG7r+VTokOqqNLWCI7OjV7g2vM
EDmxtbziHvtFzAVYUISHVGZEnGCTJ0GCSNcwtqYPk9tYcKH1mcx+YwU565BAL6TN1MAVsoHSclTl
7BDMgIqQgYGBFmxUXxMn9nuGu4Kwm0FrQ66JxNbC02AyC+LaT/2DFE4ruxXs86dzDS8PnNCemfVi
wEdXA2yBikxpm3xFVUN7YIF5yr2Tv68wImxl25OxWDD2ddl34MukY7P2DU1+xVtxu1LEen+9sXag
3O1PskqOUIbQ+PjIaIw8jGbBGWhAPUTEIQmmno1QuhICPuCY+xeTyqlP2suAFRcn401IYU7xEzzP
2ZDZvYhZevWSEk9isZ5esQRdchpru7RnTlZcgIS/l5qQqecz/ap05kpnxi8hAPS1EOXIMund/T78
9hzBD0SdepdM8I98pxQDJIk273zZfWzam6ltDBnDb4Bl6OQMP1x40CCs5t+bOvFDaLATvMqjXHwL
wz1UjkwNQXHDtOn6stgVd0uPkQ7AfzEir51bANy7+0bby0fHXd2p2yztGDcn3nQCq+8YkO5VgcnO
m+c4lfhBZe8aKI0HygS9X3diO9gfVwz6Nzv4lxZtMxC6dp8mN0CB257FKQKjCHcKQdkQVuUpPOMP
ocQOTe+LLdeuWiUECYmdRi0i0Tg4+pKAkGanaC6vQ+QyHxVf2SkGEz0S88pHYK1+PYib/srjiKOj
CSvOdnKU6LdZUGZdzV46ZD2eUErl5WjfAuv1g8AuvYN+CtIhz5SIXvMCUPvaxnG5SJdaRq8KPRjp
rpJw5V0WdlRMNdzPb12fU/G0ZnDPgXHdzSCKHPnlY1gmKGxVNN1WYwN5nXpPjS94T6UixEfK/kJB
Rmy+svB9C/DbcwsFjR3PE+LhLO2vgmnjR6UEUrlcoBjYF9gKW5vAr1u4UmWioayITP/Em4Mf+484
PpXTzy6IsagJbBDz/uVYbA6+Z6V107HrWMlJYQw32vD3cbmTOYfqljq6WO8z4PZDKk4KDqSl2qwb
3BA/l0kyJZ897e6mafkoOGNudZMLPn84qy2AR6/1Ynrlc21QgYgY44JAzsYZ1aK4W/IjAgkfbaix
hGZpIMfpsRgKnSOBJ7ZKdSLDFR2qSVTBn3vIiaUk19b5R/fEMnje2USby7M7UQBYRDEs+c+vlcXl
TY2XGTIOrJpos1FWy8+IanJISiUHJHwPjwGYJByPNVBT7Ys7rXHvoCrdecxl3Bfo74BEC9hmCV6p
wfC63hcfqHsMhrZ9Nkc73knQloze2V4eSkYfPbcVBzW/VsUBz/0TjPF6ZMcnONYDUZ6Zqhq0Or1r
zC0omlDLCwDi48icuzgRr6cEojIgZVKitvDKVk0kVW/kNUzIw9JmRRe453XD4lXB50lXuz/3ikCz
3fTeekl7206iY143564KMUz8Z7Ux7uTW/GK1FdXjUc1ZCGkZWZoKLbxX3C/EF8KpDJEnGWLBwQkO
47ftmYVWwdBdQu6L82YGHoC73x/s8V3fyktjY9kP9nj8TBHULdpnvrwWKUSxMsvx+SeOsemYwax4
n8R+oMTEnYnGHpARsqSRXjz62r5Ldf9t+i2d6RWukA/ZgJ80rESU8Ci+hEKCXGuTOMxdyJZj4wB4
ECgOyjNiN9bp8ErgKCy7ujSd1QR0CZdlh1bPch7UOHLM31ZIJ5Z4ExK0dNVjuYqNrUhNsV95y5+E
5JL+qV3yXG6ve9bjvkFHUT7Lqb8XgSQJw2CRCGrKUb4OJYFoRrEJiKyRapq1G7BktKBg3hO8BY/Y
TTR29AYYrXmKW1ij1K+BkVCthGMj1vcP/ZAotUdlaLWVlFypGXUMCj0mr7jPThI7YjQcXJd1xd9f
qoqskgXXPctJyA+pZs2bpKlY8A6huL5t/YoqRHm7tXwGuo9MMjOAmktcrbb5bC+niWizOBHLT5JS
/brdiwqtt2Qq9X7z6lMcvh7nUi8TEzWAKXvkaLx4Fz72MBtnXfAHkpROrWb0D6BFaaPZN81uNM/5
ejoGHctax8sjqCtXf+pvEm2IlldW1/JxasBkEpcBnNDYJePuq4B0ohboedDhO6mWsodzh+hW2uGM
/c6avBiq142H4C67RWEWixx1/sTUfL3kjSs04pbSZti8lgfbeNjPo37Bqr1NeSH9b7bzIB154o/I
t1aiihDJGrjrWLLsJ/HKz6pArMnEP2eQcG7gF7A+fmVUsNWJPglXby3TFG3gAeOAjMtpGWyud8NF
OUUSnwCHX5yKBlrklLKJQCH/s+wK3t8hyPIxKeBhga+QYT/39nU0AJ6UFYHeT8f/Ezrf7q1hG2rL
eQS82TbHOfnOdBIwz1TsEmV3s1HoAHOfo28DNfhp9NVxcUCc5SiQBOXfshm9TPMsUwIvXTYQqRyx
X4PANOwbqE24BszqJMd5eFc3paTDDnRVyJ0diDM1fdXrZrrUciIX/nco7HZbCPkDHwwIBxaSO9M5
Xw92LPwE7arm8R/ufyIb+HR5AeuvdqTNYYDXga6TxLQebyl+de7oTgxFx0gg275RIU+S+FhugApC
db4Bx3xpxY7Tug+Vlf0kCDbIr6viJPl5mpd3YKg+ut6yRg8nIlUt5mDPxI0VemyII/D/TH8ioMRZ
vJ1BDIMHeW5hJ/O0vDWwCPocLwocCzFhlEkDYoqG3zyYt6HE2CSJgmmNWnxMmSsigvosC/udRXGt
LQTYWSnlxQ/W7UQeFVysZetvcMy5yLYGf7cxedsjZBa6V+0mzFOVNYKu4QbLsIRpmu05tpq07v+9
lysDMfxvr6Ab4fiBkQ7sHvNDSjcHwDQESZHAp+QwpFxp4cdJ92xIQ0faWRcLqAop9ytkBRZUaf8K
MhlzE1SwDX+ZPGIBjziZXXySKapVvLdu4Ppw5/8QKGoz7l6Mm+gtyfbmSwGve7SaazbO6KiVl1wk
3wFHkWt+N2FNiczxDI1INn3X8YkiesY0zUNjBziwWZ1/BhYTBTO3Tt0J++AErWaZ7pH2O9SZFdi8
8m3KeepCyQff3ATovGZmy3cxN0ErnVE09YTfLx63v72I5IVmhyHVrKRUXJJ6sFJN2L5K+wcMlieK
tGNl3WFY0xMzhGLZRB6zr75DTMrKXhdH8khV0m6Zxs1gMNza0cUsvjoTQowEunep595pw/hUFOb0
/UuQGGPJvfrU3+gO28Wa1puR8Uf0tl4brAS+kE3WbUvx1A1eZYo6AF3hZB7/5T11mloBn8sPUV4s
4bl0JVWg7OZmt4sqgesLdYIS4zEGzPc2fj8Wg6EGO2lYVUQf0xFOZjhm0OPyGrKx9yMxdJ3xj/Y2
HHh+0uyWKAwroiCnzgPSiq+2p8U9awjYNuOUaePSIIwKbH9bCJEXVXSqa8cYhR80gt991j4or6XQ
X3a7qAX+nZ8Li3umIG1vybXCSRU5z/FVcnBwFaJBYlvQwutNfMYM1AvAX3OLNdgcLxYmNxFaTa/O
5A5L+QMMsyjtejitkFHVlnECqmue8v5N0jnXY76/sGAA6b/jTggO2Rd7uomjgneUX3XjFIW2IZKo
eUAj8KiqbUa4GeF/IVHSvyF6OP2BW7+sieRXzCfyHx1kt9BNEIAZiuN0Q4Z51PROrvSbKvv98mEV
JjlAAVvUo7A8pI2RBl/d7DsSST2W4oYyWNdEE0Pci+cIbcRfcKXJBQ2T8dXLwcpCK500e1CkJSue
Wpud2hOgHNMyrM7XVVrc3jmD3D6i2U/lh1deB6jgrnLPvBJn2kHfybEYb35jynURTqrpMRsbCNaJ
n4AQkzMCvPLaau+N4b68qpmLFySbekZcSIC0Ssa9CTKRsSecl1tW03sxeJH6mEJI9AdYgOOvlh6q
vH2HkWgKi3avuUM0yxVV1eQHfC/k/fcJkzBRbYUwag77V8mmMTqrWURh297ztqODqoLRya8wgJWW
3H03vVzR8S2/uwbzMBBncG5owASos9dnxPc7otEkEmTSeySFPjF7CKyrYJu7pdo2g3g6udHHmSkp
3WEM6RwugFxCB69zunNt/wdmJxYwufJ9E9sG/YoCMq6iKFiWUtWI1gqJLtvDc0ktK7mjjLKpjRhL
RcnOQO7ImAo53PiZ78FSu9zl5Po5oipIOv1JdHswT1XfdU5uA7PpkQY1pWApXHkVTU2d2ZZjQVnl
NT7zne04w8YPvkKxVJqFpneWQyKu60fg/K3gYKeUKpVbocz5tJM678uZEidaSOZJ8ubL4oLxpaQG
ddwisHTQ/rbyC2u29beWww6c2rSJ/SR/3w9UpGEUWTRVqsTQtXy0fkmG77OoCfVRjYZnl7G/9RpY
7rCnJGBYTvCEOm8Lc7u/DbP6leuPdD7oVmlvEn6QT6GWWyEtPbXex6Ncnx7fK0xd4xjTgfUAaWDR
TFpfHdluPHtwAKAJ1hNaBNuW4jaEGWy6st75DKyQZlepLRPxCK9kOhcamwArGvCelfNR5lI5SPF9
d+STNZ9WAMvv3Gc/Q9sU4F1o2eJW30/ch4NNTFSOayPKKpTDZz2D4F2NX2Ci6JI1Q2+Y8u24cVlC
lPb0QKK/TFRTDTPkwNGfWPLck5zhlulM//axbxj2RT3mGguEbVunsFXZRDfOpMWtPB/FBGowGIkz
VpT8cVGlmcsj26hTkI75Oza6zIlgy+BbG49SPaUP47zKwcOeIhZRflyUSexFCvm25Jp1/ABIEux1
8oaZcyCIq0c42N3yKTDgUKtDq8Gvow4N7e1WW4VMWiRlqqXH0x7lUxwOSNn/N1mquht5rn2G94de
cfCAFdgMUZslnc4yxFSEHLRMh2aC2YOsPfubQ31iNmQVZD09EFnCTlofJQtUcq4u4UZNnJ+1HkYl
c0gKFp113xLtkd6VYaw8knwdaibNAP1QDxu7yqLhJtRTruJ2ac9KJkAf5muiFnP+F2AI0IU+UrW8
HJF5xedDSzVTO45w8zs/4ckm97/WCgngWLmlmOH8VOL1PYYVc7mhwCjxDIYptHQPWYas2twH//bn
HPRo7JOGPRgwHNh1/iagzQ80MVQ12HqyNzAZZ/cYmTB91EZKwdZmXZ4xrFT6qrknLf5HIQoOzkqZ
xP5Mgdfrp9zgg5z1DTObNaE6wvGC9o47ke7wUc/fVxjGEM2EVfbzCgZZsGAcu6tY7IfS3V+6mhCL
ofYwiqA7dcoRACh5qRKBkbPn6loxbTOb3tNw5kgClphgKx2zstzc254mgWJcpjWZwFpQCziDgVau
bq0pNWNz8Oja3gaqFCBWo2d1rTZAcKbY3plsGQ/5SKnvZZifV1BM6Z/ZikVqeFteTp4KKkavXck/
C9R+PsapTDv9XASBfuZ1ThcYLiK5IiDWM9zVrIpHMJjWldp5FXArrSEIjfbiYcs9A/zFKMtosEwK
KkOFxp8PB6ZaWvitZzuUJ4K7BbHxFUKjV3LlcKzpjAivMg/ADg68KchqMDXvYSt+qFKsYFLfSsFn
ZOo4XWsVd9kTuAoPGFKrtIte14Shatm8BGrS7D+f+rgmPB7JDwwlc9qRu956YouM+e0Pfg3pHorK
e6co+6WYKQRWc14aSvbnUtoXYmd6c4L3+DMlPI/u1BhruIedVX0XTufu/tSKBpicDDuSxQXX+eo4
5VAxI+mw7HBlhoWN3RpXhVTmQnLX8xPzliALevy57y1Dm+CtkArxJ1v8bC4n2zEpparuSGSa4aYx
TlQlK9+VHVKKshkZbAVrf1bLqx4jndEccFOsKBrdlWHjAf+QcketCBJin+zp7ZAGhr95NzzV0ZpN
7hnW+2vw8oMaHJKJkIpQ9ndXGJ/prlYgR/uQ24elSzfPIcGXFlIxvbQRDP+XEZUesFxEhk9ur4EQ
rfFvwhIQbYViU1xwmZIE5JWP/CcOg/6wpgMh+cN01VNElLxL5f3O+kYTS5lT/9YWrh5D0tJ+ALfa
kGBhvR5KEPSsa0FViljosFzRYEp+7MIUBhA5DNiNht9sT6jfOHyR9H95qNA7PLqoqsFpDGXTdcIA
zPJ6HoC2fD/bMJD2eznVyTqM/DxMpFFg0lVC2lGdLDIwqAZ9MbOkmpSKU0vsHlT03ufXOwF4TzV8
8fL3WyOcBXlewommdq4DYZVSO/ib2nNJHgtHqIAZRdD0VmVUPauFw+U9x2elJ07e15kgd71rKh2f
ccIi0yXF7Eab4/d3xdiA6JFsbXOl0JIe1QrRa6QWX9U/7ElmWQDonz1zAalyBBNinHKKACMe15VG
fRp+KefRczODSbzv11dB5kWfJ//LeMpFrt9t5pP2f1ZX3GC8hAo3Vx8Q9SvPH7BwE/WRTWpqBrJE
60sZTbNxE8PmKblZfANuCy78vg3E+UgyV50tf2/gX0+N4H7fl1HJgjXjEaP/uNDKEMwYbEg83L/l
Wdvo4ucz+vZwhsz9ayaMXl5HdZcZKBjz4N00c+YoQ/209QPeOoBkRNNkPUte5jBy2cM5qvV9I+Tg
7SujqCYxUc+RBPrvsnSaX8wAghtDbnhmeKsYNeMfjUxcpVvx7+VStsT7ZlxDpW3kSwApoAg8MP2B
lxQXDOYeQsOwQULR4EDhP1NIx56WMSQOJ/6wUIjJAWKvwYmzfy6CrfDHOvfrYzi4cVHLoUphtYLb
G8THdjmmrXdIHQARikjB2jwjN+4LHICLnX09EwJEv274mKxiC4K3ukuhVASWN/bWOLIP5/7q8MNQ
E3LrM9+HPfFCjIPjeLh6B42WW5CWdidDY2MmNw4ufuJmY87lfGriuqAgcHQJTt1Ft/dksk6PuQ/g
iGrGvHzIuUFZGVeGyUexhtAuJ+y3vj9qjhlmwK1pM9aZrNkui79GpAOGPIQ1T8GlI+UgNl5sqQFQ
wpA4gGawK6+oXxupr8VtAoHuv+IcwWsRYnfMmRL8LeEyk7AfXdG8MY+ysbGCUOf3sAOCNCbfcaqA
CxNY5Jg1UEx7NJ7qUBnZWFOB3k0RVHb0PtVz+CKaIsD/MQrcFkByErr40eSRp0NUi3O7qvShhRhF
uHxpxLEOH/V8eu6FYjuUy8gIJDkeilTvefWa9tJRTFOar3qlCTJuvm933hh4aAQ4dB+vqmMiuFNG
NsGThyC9fdh5LZhRTMFA+KP8ua8MWn9pHpgPvzz6QDDcsnV1DcSrVVWR+4g0ekdP7L0QHQRNtoNT
pgfHLdWrscgZ9C9a1deOJnZ+Ld0WWucPnOKkC0Jim7x3xb8O0eYXFMxvTsHXwZy3g3jXpwCfNAwU
/EeUXEwRKCIW7zkd5guIq6pzd1q+7889SEtK03MLPLRKUCxOS6oFD5rIJuhecGaRUNU3WRukjBQS
MaixWWXbdRU+b1XuWvawi6RjrBbYgpjVtWL5xMI0RkkhCZ2mprRrkXm+Wuw+qSREiqEUT53y5K4u
lA0B5i6oCDOElMudLjmYW93IvxgqVKTr0uTVGMZCaFKL7el/S+Adui/+z+k4soXlpqlsM2qDGsim
P3gcvCfq6R92p7Fkl4vc/BhINEDdYr7nTG8G1fuJA9HhSpBjYZFahBXXXMBxZYOwk6VirW/QxiWO
tleHMBZICwwE1upDo0mwRprY4NPVA4iMCyWfzIH+w7nZXln0t8CAU4SCbNwioVwM5M0Vz7z5VvdH
rE+QQgOdNzwf7HJPvuXp/XIOvZIhVUVUOXjYor5e8hlM/xm/Dzx4TCPtp9RYjRIfy1SChuH3iYCf
Tx98YWUrc2kpFQ8NJAAppwX9PSGpzOmyMwXgDVVup9Kdx6Q2236RIKLHbu49/VeK2Qvkgp9XPiL9
14PgIm0uMSweRCqRMcJRUY0Q0/64TqeAYbFh067B0tIEn+SbgmXFtRvZkLPy932EnNRZ8olqSkoE
yqsEJQnbSZU8D0uXBEWpGwPyKr35/QJDt8bSGEmC9s83X2czJv5FGmzL+Tx+qx13Fs2DbXMNurpj
Ogulc7Js5L7XV+/1VqFw+xRan84BkTRuVAyGJ1lihDFvUWIwlHiwPJZUqQ0heYe8KXsojo20eQmZ
cCXkdMXA2PvYu/Dyng7ao1VIDB8CMixnEnlIQa7Ot0gwK0XIeWs5FClxJLBb1TVaTSygcuojrr28
r2xYgFjhKbaLqu+ZeRf8DUcsOgXg5YCkOSRHVWtPN1DCN+klZSK46D44EvrpHUTUTJZSwZ7jRJdP
rlFLSkQEh98ugGgLu0FQEZIGLS5eC1Dj27koTzBsxwrumHjBy7wrwQMmyXQlnqL3no2bcuS0gY4v
Hf+CKDkUXcYfYRl0YjMk7sbdmtue9uadklcN/buIwP1TrMBASgNXRRBHiBXS1wdH1rITc2FR6piX
z+LdpbYVrdE8FjQKhYJF66oTvzTmBVQX4VjK81IMcc0RKJaoN4FlpjYwDA42cpSLad5oBzY1Y8Ji
9zCoB2wyxd5e6e1ytVM27km8Fyiy08fXm+KCQpjJnxc006k17sqAvTXzoeSdywuXmH41N2yLYvSz
1uB6tD0V90tKVgFKPyF0E/sVt0cKRebNDniOWAEhn6GoFo7Pe2phVlRgru094qJOFuOGRwKzOgk7
HB41UaDT7PbFAp8RjgUE0bWOni9/Ge7DUYBxoEEEGpxNcAL1yadxyhptEkV9Y8egis3dDVFdnpjx
bRUK6hFlPBWNVQ4AMXAT0ZCzzhnFcc0RzS4/206IDvdCxyt5gfb4od8XpcVJPqP4s3wsDa9GWWEw
EKfnkUOapoM1ztWPSZNFNPOes/Ha9pGAysB6Ra8XYMEfKKoi9qXNfuv8l8l3JIWvrOHc6U1K4WH/
uhje/8DGWDqcpSyxFrAxTpUxfEOoZMboocJNrVrTMUCWS/OsvF5/37AycqirLea9Yq3lGM0iQx6E
/0J5OPya66uxdDmoC7oKM1yYXqDjMBs3f3k7UsuwwroyxNJDs9lKMdK1ziy+1b0jinhxgcfQlCND
uWbvbe/+D2Gf5R5EQMwesLFKTAZTlWwFDlrM/qP9eB00KcYL7POwtmWG9XYaJrXpkammHI2pVsGq
Kebqlpo+uLZBhwIn8RrJID0dix+96HccuAz5gdw2mUKqXEDr5sB/o1dyJ6mGoBq9eKH7wzLmOaQI
utIe1HLok22SQnCqy75fw3jr2lhEQOEeyL35Ivwn4tRGP/boMLuK8bO/9IhsOB03CZCNvJk9Z86k
tQRzozHiuObgtFmL5hmhKT5CgMB21+VCQsD9LIxUNbuKvV6bZrFcJ8kbbwRNb6o4KZ8uyARg5arw
0Xxm81HjHt3nyuUwQt+FusDpjTwogR67nY1mkXqpxMixGANWIBl5BGu9Nhf8lWQb51/I/sKjZh1U
lLOzgiRXtwwxIk1xqg60Zo3qIKeZR+PaZDZW+Z3339uuq4FJ/5CiTyQchrXPBWd9luediX6bOgGC
E5d5cPMsr+nwN0nkwTDOBVJdz5CzugWJ5ETnlAj8yE/Xq37YRfWsGGRZIUkDE2nDnnVnVO6NRMjz
kdXAGG4BX21AovxwvgYqRO2jsFNceRj8DVOTSA8sySBrzSJjz31lj9/iePKv8fuOl7nrOFfwr1aE
zYcDXnUAO7BodaHXbJT1PgCQsCttHQJRgX4J/FAZPHnBGius/U46FiUtociG10GtW238eJv77B+e
0IsKeeGfN7X04f8dVRmaQmMtpXm5212wB3/EBraUlOThTygrRJD80Ywf/OR/zNWhkU6fH65ytsLT
JiUS/UZzRvojzOZLFJHrxtAIhg/G5GaBvKaruYoT7mFpcM5EJg6bpjLt264PjZfu+w0cFRQN5W3b
XOQaWPKrIyuqIrRmMYEceEip7Vmj/o7P4u4iEI7NZRWH8BoaeJcdFUpHcrCk4UmLwrfV7aWv44te
Aj8kHUpuQoX8LjCuxAN1pt6NRNgIa3ug7f6R9g/8wr0ViUsw5r1lCvHjsk9bAtKRB4Hjj/P14DIc
POS0mF5Y9d7RFqdk/561g7Mqeb6E14NZMQG+q7mN5No5K5uP5t2L1Aq85xcVhH7J5yjs43r4pmw3
12NWJ1LggTGRwKKakgY0mz7zuoxXgNLJhiPDs40GDCpO892bURl0uikGtQ1eP+7K9BtUCDguaWPq
MjF3eToSL+MQYqKCRHv9gJ/qBMqOOYUEXhWgNy7ql+NBXc63orlqImsGAj/6WABU6q2Vn/IsFQrC
/fwo0ym5p78MxKp0IuRfcCMwI2WikTwEaqYzF/wY07+PeOUu4ogTuQM4K2nmZaTvBNfmXW2/ynQp
yMfiThcUfMKULj06ZeQz/smKchIKInD+EOVEp4v88JDrQqbDtneEcq9lo5NkwjpSjeknWtJ2ntVM
os6OtOtqvBgb/B8IBrvF8jCpisz689vW7TNJ6Jq3DNraAm9oGiOZynPcQe54FaDM9taQlQGHzIOz
DgHwwoEd3ulytvJTBicyoOgHml7U1SwqBhm04Y8qIsunRurEFRYME/M8iSCVquEdYXLkJNCqpzlR
ae4IyW3j46rFjV9nnvEotxtVlYfE3Gl1mOTRNkWL55Tn1+FriIjeTK8Sxaq/0eH20y05vvvM4lJp
7Soe59yJu8hDitnWhpuJ2MDE6aLTGITGSeBkb6vWj0W/AKFVwV4/iPQDKabUDuP3Dm07r10FnW29
Tue6f5Ef9Nn+Knc1JjfT/rL0FFNL0E+/guFL/8efxSHwvI7FF0yZowledpXrBQNv/CTTB9GWm257
5SXfc3fu6+Wkp3I54Tk3bgiT7wiBLy2Hd3atUrW/iKLs91vR3S838oqg+VEfPRofwpFM8QsvJ6RL
v+Qq69wmVubORLToOJYeQSyUsuaCX+Fxhv1J5oeeTfR0ou6EU9jhkxh/qpGhQSdbei02XJCXiTDe
4ZNkh8U5C7bbEejFlQRE2YfP3X/MEqVJbjy1q1tOkwwrAZU03F0K3Z3RtpRYo+h/RAgtdxEFr7d/
FUmsy0cEWeAhiPgwqAfV6V2HUqsbomf17Et7fw+FkLge0PO9qFxBKxk6mplEbwFf/LNtBiTWoQrQ
V/MQ/d9UQxJ//jAnARFPckEO+jIj/BALk12cnwa7yVl5nNl2ZPf55SCjZL/rtbuZf8y/nvB7t58z
IsjycCxPJyOVXbl9hkz9YHDzvXQc2IdEyb3OrqnkF9IxQFi3KmCmzhd5Rf9nXdXEwfpclduu5uQ3
/7Dzs4+vfzX2GE22EmRBbFVf4APTL3wQFKjMYATfWkMZDFILWcTweeivNtmNTIYOVf+U6tOTq/O3
9KJ2aplTlcFLZP+lWtJXXW/TzoHHGtoyzz42pzj9Kdo2Drdxla6/uKM2gtJ3e6FOU/ENnPF6tbe2
U+bu9zyHMMURGZ/EQ0WdHVvr2/SA1WS8A6uH6SNRm8u5HyXe++X81yLNk3OGcIP5tpeW4/jxL5gs
LM5Jz9G8LOBA9o92VhFvpsYg7514/Rl/sMFIrS7KGeU1Ta/NI4aQf5SDNyoKi7EdW2SymS1ofSp6
ZBv7st/2hAhuL5W4DpJqCvUZI89ZNsSJIy1eWLAuBLKDqFVP9CUs+XpxmEGJYgwoeC+EFTKNu2lf
7LZjGx5cZRhnjb6h8uyr2xja3UmjB15uijuz2mpZaQ8/BsCZ6gIgn7cWIjCg/+hku0plxJ4G0plG
VlyWW0+K4Y14afy2IVf4BSVz43kzWMgIO28/oo3raEU3aEKrINqie1xBNlEbXLG1GNLS5Gd8v+nl
w4Hh3X7/UZyQbMVjMeTxHrFWgOL8Fv5qjiKt7q7Q+m6SUacWEK1OQJzgeZQYY/biSJnjyT51o6if
jMPWkqAUSBTA5Z3plFUq0NlK6yun4jS8vU5mXQftXqEiwDnMdbtSmOwisL6yFCalQ4nJYAA7duOP
TwvXeQnkLWJ1Muc6IWTBkuWRsWo+4GTKl1ItT5IZ9VDWvBuLeZvZCor4xOJQJEqpQUsTKnjnYXn4
4vLlBTAh/b2PuYFq9yiid5P650cDz+6CpcKRVrvwREv5W3orwvsP/ex/V/eZ2Zgs6v7A5Y16i1y8
uC5SvAHyzvGKhB+1xJnb9alJOJRscuP0GwM4LmvEuTPmlfgJi+n48wB3PwFui+yJdXC+Ru4oaf85
Z4jJs8fZQPCQ3CAncJ9EPnHNjF3DghMB5UEB0Cw6X37BKAlmjdG0SGeRxrGvVPlZ3Au3XnkMStDi
jq6TvDBwYwV8e+nd9pY2dtKctgk0E+cFq4EK4fTjDrqy6Mzyil7v5x66qiZm+QqQas2srPc2T4nn
XZjJysSCyuAaOOf/NuZr4b3EoHMkX1n7EK8e+W8i5Ct2M2Yy2Nc9qy2mT3nH0HXavHy3ep8IOpTt
VADa0VqbnnXN9SjvG5XTjC1nFnDk0R12pv5+wxrL/tLrMxY/bPILuY7VWNskTpAud9MrlC0TBMqB
zKnHl50xDAg/CCY8lLhSNAbIFBFOoNA48Tv0rVhPpyB0mH8nLyu/1AZLCNxwTBBGJsPkgwrpX/k0
x1ASXxWGvj164YlsEPIzW85GhQqp5ND07HS9LhG/2GKhWLcESxjrzwYDVO0lwpCR5hzOEBcm7i4K
PgXN58tmKQgF5uISE/4YzSTiKZoCkynqPzCa/oHq2/LykU4kQDRZaz++Easo8dKKflun3KUgS55k
yWG8Jux61n7s9n0GymDMLvx39X5cinSToPVeI61tFV9VrufNPDGWOMM0hmenbEfCiwz//Gd0jCbv
sIv1HIiveaMvJ0ebnu5SOkZKWqZYX1a8tlFNlTJT0s+x4pDaDh24VmvesV8sIefFp1lAXtJkpHTG
dmUfuelaSyjPsF++GmcXZVJ0/2rj0hIQVFlBV2JgTatdAv/vRKbd2wIJ2rHJriZj7UEd0t7yX6X6
C2nuTHsA7TytTd2jmtF48Craxo2C3/Loz3qnlnBF7pZ/enyFjYU5D/10OpLTG/d3Jzoc7hd6BWbk
ZMa51zfPBruXTzZxUZJYuI/EhjYDPqAmsw0eC79QjnZBh000nywZqlzzesGCR3J2sesHLXeVEuFS
pJSR7q0OYLjVd5Ekn3B/mlNKsbunZAX52MV7KITX7C6K2HeI8bCwzNRL7f9vbZ13uLDzizCjI44O
OvC6vWQpXoCDiT5Z6DT0SU0qbl2R9NfQtz1nMEMm710YYgf9uhZU39wZf0kC7CVyMkZuLJbgbZq6
PUM196ukF9Gbey80sw9UL1tO8t/mhmw7zY+LhLKmjdtIO/0cZxcLg2ofPKAt1VEYH7abdZgSift4
+zuxkoKkMwGHbdc28r3aRkDCvv46vGazIg/pkx89H2BAn7ecr893H4GbCDcmvuMJ+xSli922cX/E
eWeVUCmKRg40gneq4H9vW2mJoURH3uhJHkh3kQRTakQUMB9eArkqzrpVYTOzjAmAyQheIHzgagZl
d26bgqmUm6+/8r4ATZyVTfngmuLpOspYhkotMqPY9EvxqjLGNYiSYGPaCAiH+FGeJp2afCS2jwv3
DH3gDWSl7uVgNBKyxT8DpF3ID0uZV1KYH8PJBakpGNI+oLvm0k8/L2EuEGsMWvfdbRPcVslJK2ZX
3QqGc6BTA7rUige96kSwfDMjqVF8YkQh85VQ5Muk/hCJQ9Nl6Jxt7Yhztg7/dyogOPUgbcGI9t7J
uyVg8N2IcIGr4OFQWZ3ESwwx+70ytVCUjwGn0W6osH3AY4ZAMopQC14X+aiseSpEop+KOEU1BVHD
MBPEYCxcpkPtFQ2dpf7m33E8sVfIdTsemloS4u5juokYHU9Rsmb7w8kXaeRNtgH9o4vRZeFC53bP
C/3dalDxA75Hv0aCAnwcn7z7MdbjDn58HGJ++R7ze35K1BJaaQ4xO1PdSGWR1LUD1iu+9ykHv/H/
soBYsg8EZkYRMvRMuiB0w06U2WmJ6g1AsJEN9b65VAGHahVMxKeMBHbed4gPCZonzRJ9S+yEu2bo
knUqO+RaRhAGNmvOfo6CMeVZB3Cuqfd6Ytfy3AX4qnxm+a6H4nx7db9aJUEa+Vz1nZX/znX58JJj
xq7rFhAZgko99g0Vs+CNDHDcXbmcoMQSE2HarDVcImERX0tWW3/4T1s11QE93Oa+KPXnwmN5mVq4
lEiI29pBHWQA/MOh77PqnrNArbxvX8c9lOyM179Rydx4GsX74LL4WpI1vzb3FD3uL553QeaNKil2
Br+/IPtw3/RMbVfWL4CZqwGJ1Askr0niN/2haX+Tn7iWzme30pzPRgeOb6MHZU0fft0LXW1A7ZFf
V19afq4a7w9wdK83jdTh3EjeFtB3butsEVutSUSdw69Ryxg35bdRmiE5/fABDUePXiDbddwk8YiE
Q6adsLKNR+LUV0ID3XJT5UBxLDROvJWOEaVH8aMHpXmV6G3tPnf11w5qeXbMhB0Daw590JRNC5sd
czRX27mxJW4XvNt6HlFqFZVi6ilRQsx8kRvC3SCGMl2MPNOJJ5KzyHCDfqSfczVkfV+kMyu69uHm
IAuJkTz8yqJORBzE0FQPKPvvzN7tD8ISfgd+MN5q+dJfmQr3mEnXPvxlSQGGUlKy+pppetLnm0Aq
C1/QMAnK9btV/R4U9KPRmvK31fIe6r2s8xp4nviSLiu44RVZ1pwzIqxT41pHkhWt6gbId7XrgV7i
o8lbYECke4pcJwkOlr02cZ54haeDbsWbuRTrQtXxHYFGHAu45AfYzhsDgZAsxKcbgKiNcjidoKfw
p1cTXd4UiNKbpQBfBWl3cjYZX7uWPwhHUTS/uRDgs8tKNZOo8d316N0G2OkZ5YkyOdzexcTmsUch
ZrhLWqd2RGTzFIT7lSESfBQhI1y62sxF0JHZj/LtScBBRHNRWUMPY7ds7pOXRLkeftSClbL3/pBA
Aga3rI/5h/2aHDv2/IbfcfmApR8y7VS89qLOmIbX5220bOnOa/uBOjp4c05m49zfNDGJ3eQzU4oZ
6nVErUh8LrE7gGur7WmmPFTnot4qus/B2u/qsGd4Bi6f+Jfuptwg29jZrQBqNQxD2Ba000AnA1rq
tonuOoWIFlhtEXpEjvGykL25zuYwr/bWIu1pXfy4h4dJ+dbrB+s7avolvlL9HZo6peQtA/dWQsNl
5AnbQ9qFOl4N8Iv7XnkjFpyiYwwV5NA8azcG7fNL4pU9tsmV4LnuVEU++Zv+8Gd2BdTBTq34PZVH
M0GD3CNUJjVnswTadZClECMVFDxkGcMsXCcSVMMfijb3URLfFYx58ZMQTIEt9T2sOkYkWW4WiEWL
jLRF+PjGzVtpc9ycfA6pPQI7PdEaqsBgndpvQiv6FZX3HN4niiS2cqbzm5akwyVV8x5UQ7FiUpBA
xREYwCk6u7TqLgvdv0CT1ffGND2gEv9O6j/9jPqbqFaF8JkZ4rSrVQ/JTNasWePR8eM/c/7vaqRr
J44KQfGmJ0s0NLfm39Ln3o1hvI5Puhq/CgX0Vwc7vaKcfoQr2Rie/m8uULiWL7CNx5dzFXJw/NTw
CxeZABQ/CHydv9xRI5zX0a+HZgFbMKt1XZufirPKpjOMv4maYydCZ+4SXOaeV571rm9yKH0bfbw0
/24qiMsrei6pTnJlL2umPAncbyczu4JQzX0ca1RUb7/S5XAJytv/Xfe4YbIuNjOi4GCW4PbLl55Z
teJauqjVWJCUjuxTsFW5bDtsSakO12tXD6D9m1dGjTQZ/iIFRbDhVJLKUGdDbANtboUw7U3+dIyJ
a9wmlrdtPk4egUawSFs1dg34txPWK8T5hP8GKFrU3ixbYE2fw45MQp2uWwx4hnE09zZrkoQ27Yw5
1ACpxjRYDhrSGJUKWZYstmC7C84oY9Wh1RnVC9JhyB0MS3TUq/Z9lLnfVd0QGfqzha36QeIJDyS6
omY43RSSt9AmGIO4FchCRINr6ai+Qt8qjz8PBvBuGwMh6bqxx+LvsuSo5nyQ35j+3N7WguKiNlkq
e8lyrbiezEJCRZvwNAt1IxkV4+FfeYQynGXpBnvHzXu7232Z+fZrJIiboXZC6j0TyEH9QaKjFNU5
fq2waG2sANPBqUlDs/G7L7CBFXt+4iItnHLsj89XwD/B9AELk12XHd6nJY0ogLLiXxD3AjcHPGAu
q7CszglrzLzjnjB2/sEpIPGSNOiGyV/Qcdh7iE13RSRhsFhkdKtuJNUlOp4G9Hzu2n9dgXgPlVnH
THzxmchEocDE3jSfKMT9K3KB8HivzklVuNR0cnltp8T20hQkYmKBcEpEbV5R1P4unayFg8o3CjZl
aKkI7CUnNAHhqYIgVH7xqpeVoVVfYpCgmV+wg32uHbQlnfcy4ygfegvbSyqWs908gDQvEn/JJcY1
kkKepQK8CUi7+aRbw4J3cwntrFzMiGHa2h9gISNIMugiQ8J7If0WDhp59eQ1JnbS5hRDSv02gPLK
8PR1FWpCrjCegt0uIgFkl0SapJC6Ip1tWoI0pZeuOAVGommYWIh/dq9iMokIUJUHF00YrqDlMbgP
OlFe0JNt/+f8pyGQPoRBQK4vKR+cD/AJGRDajkX7wQpj+2oEWxrHW0F7MqKzRx7tcUEwR/Y/eDl9
wAuK5qkEjnXul79E35T01MKjSdU5tf7p39axr6e+iI3eYomkImiGzN7XtOjurG3vXsvTTZouQtIx
AN/nexy359TiZJBT0xc/fO5QJFXSMtRqPq9qK7K3T2obYUQgd8CLYhonvccpuasKxF9xiiRxeO/n
uunVA+DUTVQiGojmaXmcAJshmU3E5j9HmjKs7e/zQflTpV8KFjoahpabigHcym8lazxOl2neMByW
ogVmniAYByAexLjHV0q0NKqrFxvga7TAjwd3JFhREZevSU1sDXPap5AubWIIoJiENjF1YbJUp/Ko
N+VRv8tlQ2JhrCwOHRyj/NpuQV9UinvEA9QeMeS29mc8pNovY/v0hbVeus/rRC5LY2kwQM5qEgTj
m+5xk0ny/k933LZ9iS80DVbXzyWer7uzgAajTY+7OmHyZ+vBGt2PhnWGWmprIJn/EvgEVV3gYTMJ
G4f9zjdKV4D4kMYfXT5LiT1axagkHcYHwOyCSwo3GMg7v8EeLjB2E0cVMTGY7XSZ1VHlsd02IrLH
xAGrXmgQQWbYfd4hiYlANvxJDRMDxX4vYdwvYDdAYN7oDT/M+gZU0UN+tB5ie3STfb4GXyCJm5xJ
weJ4mtGary54QLjLxci/Gt0gz4E/3JOLPOcB7wi7w4wZLZGV+/w6JWAaefz98GLi2m8s1IFPLuso
tA0tVK28agvthjDeeNLBY67CBZn9cegbvxibLoikne86NyBN+bylL7h5TBef+Y+EwJQGZ0QDm1Xt
MFkiYo2UaS9AsauGGpOgsbWxsy+/fwu076iPllv0r7FCEdB4Gm3wXCxjDShwpuCxNOWnnlBGaejR
193e8pxV63X96xR0b2bBg5o8rp3ckGhB2intvkztLKp5QZxqznpj0h+KkqoUazdK9+1OMcllO31c
+bov0onDCkpJ5TcJoGWxGjdlBI0NPhTz1nvW4BRCZiWEcFKp3SF+XgfYG4svhJLbN1yGs5NRcdDM
d/bWDSc4RtRVrKLwMZI/+F1T2/xjN/xntds5pTrC91yabJQ0qHk5fEDXb070kNgiEZ+O9bxBqWZt
578VTUs4oOm2Yu6RpNKibdjvTlKTiMQNYd6sqm2s1sHeZOdx5yE7WDcUoqCWJTPaCil7KVLUbPEl
2HHvd10bJsU66vzOBh9ZeoHz5cEX2MYMvh4e4Ef8CX9R3S43lqkl2a3OvrqeweM5oblfnRF0OdnP
caZG3Gn5UHfND0HE+jjrVdJDZIehzmVs2bh5xH1Fv2XqWXnKX8RzMQxPBBlI5k0x1Ttv16+FRAND
ZzgdDl5HGSy4Ib/GDaTvqXbm0z1nagDc0EqdCQXYy9I9KK7lR0OA8Tmloc7bLbHvpo90XTWk1QYT
Xd4BKy+z1k3dNjPZq8/1t3S2YeOBiLdxGd8WaLH5dtG2iIxRqNTFNsg7zfOuFvhEqDxTNq4aX5uT
d+cmHGXewAbPPnmuwIwR68R5SPEhtROrwex/qruh3YsmOd4vM716c/RiQ74VXO4BN6bE9a08aSyZ
rUiuNCTTe3kH0dKxN2VODkLQYMjejJ2+ps2qGGjRK9q1fsopAA/dbv9lIUOitmfpRLq1z5kvyaTq
0JZKl8moa1qvw3fnR1+4HGFHE6sdPdaUKMTeBJRpyDFEHP648+7PBK+Tutr3jtLVrvBpkecp1Nvj
FhISGxpEDBLWEyJun8wWEloAvGtnOZ1Rxkf3fvxoni24vZlOY4Ff3gRsbASdV+SbKgPwdoHj1CwH
4k/U1aD9aD2JeftyMfubR2zkdx84U4947vDa8PKfpcxPFxl8ma7Tp9nnhbSIOD8stMybuCQ+ZIYB
KCAtBc/xAKU/WWSG32q6owWNo3NAnF9ry52vsdxGTVy6StJpOjnePcQ6D2bLxXJfT7Sqp53INxjH
RTxN39i212lSxpv6o2iLnkeOhSvSAD7QYVANtbv5VBeDJ8pT/op1h76RlWX7+x7uRw6/+pwRqV8c
OMbsq5zsLvsIdmF/5n46zMBtyOZNZQJhvBKQVmapfSrNBp7wsJcWjsbJKnKU0JD1qQwN0/gJ9lpu
B9AeUyDCGVcmTrIlWbwkV8udvP4RSczkCbki4ZFqXXv+5zWHyqHsLnq90vOV+bvTEvro3BSBO4Eb
QL2uTRujtdNC3rwtaIWEXCtJDNNckO095z5ld7cx5DNKmJSnxTCjiL3/Ab4+wULQEFvgoQtS/kG/
7jGfwvZ/ossXZaPJJg4l/c4iiIvfTgkZF2aDQu3cEH/VAf26SzKwZOkYN2KySR8Ulhw0vx6+Orbq
bDt1YCV36G+yhIFeszTNeIYap0Uagf4lbI9hBwoI+dB0SBTbejMPbzHMNfgMC+2BpyyMIo8NH8V6
VYYLbYW1fdi9yp0oGw0eUGs8rftYzmZDj7h0uaXvVUjjtnXAR/nkoXJWYj6tr2kqUIvPrP4mKtNT
2czSQ+LjkEZc30jvab8Xh/7Wn13yXVgG52BvrpGJWqncNbAetMkPMj4rfZV+OMK0xcnVWpfqWSyH
an1mducmgq5VmAYymscahxzcVvXVDUhh+dmhq/C8c/6wRwKIjtD/DzrBZ5e1XkUlsFAs6fHbh1nq
691ZY3JG86pLT9Nno9gGT/TkE809H2nj+p1VZAT3XX/3Tt0ZjxuWH+cQO7/8J4sYz7/2foI4oET2
WxF0zVNXlPUH25fnX+dlIQ9+506nyTLjI+rZ2/GdDbu6ReN0itg8Hu+fxkUpohTK22fwz3PJhN7j
xqLAbaJ4k52xwsfVO06lk56tx4jBd0tw6wrCMHZb86HX4EF5nLLjfyqcXI/H22+xSaDPXoAG/qI9
VibDnb+8YevD5sJmjo9EwnyxyMnPHPk4OreaiaJzh9C9jcK46wzUzN0HFOHNhWviLW7HW8iXlRAX
cvrKvBGSAjipxEPrfq7rA0zkMziWOVGri2g2okZEDY6/VUfDk3gE6tYm7bbgC5gBvdtJUo5eBkRn
a2Kvcex08IF+WPOYw/haU+JoZVuXWwp/H7b3Cz49ukYJGggOGG9b4Y3LKKxbtgYirHqhlm4g9wy3
mfMtQKnjk5SMtzlzMPe0U9k/V5h8KTPLOJ8EF0t8hOUcZxnHtcpsvBwPWJbj3gtsoDgoHTS842id
a7PeCnAq/7ASNQUOl4j5ju/I4tUdGRrUxWexN37NRk6JHBJSXVjl1kHxHLJuHFJ722bsPkkI/dN8
d/2msHBpdfctPLfQwX3wiop2hK4XK17zvr97z/2vzxRIdcbW+U/xd9g+mhiepX1uZ40GA2vF455E
XE3y3iev0cfD03Y4JSScLGzmpH4ir4lcSgcDd+PCr8Hp2B9f5MjIvoKDR+NUmyWoc0Quq4h/JImK
UBSEarS+rW8V4G/qo6pnNI3fclUqwRg/wJmwQliuBGZV3larB35L5wraB8c4sg1MRsFCjIFa1Bwl
UyUNOulRzBpoVaxC10P9qYv0KHHzuxl1eWAdqfI9TJaN8xdBG4gZX+z2y3UuHEEgmw5JHdegGZaL
hmuZiKpbFEUQlt8HHV5ogmR/cK7uF0gGq0N3nnpfZu8XMYgoBRV3Co9MHz59/lCnFeZjVfazz3ne
6wIg5+sTW4Sd32YThBMFx4aDpIH5tArU/LGnXMOCqAXP5eSARY8xhrBjJAugp3dfrEH0jYDAt8wD
YoFHAWRrJDAMJNkdT5fOclXEk8x3fLpZhO+jghK/TeMKDpXIs+0Hwzw2lKDV+0pUgk7g82qvd52H
5AJsnJ472ibdKYq/FO3AprhZOjTTbPJF2T0H+8DD2eyOexW7sZWLGOspXxj+mI8nT3gZvtEmeAst
TLYb00ucl9wA9yEM/KUTrj7wpjuL/+2MVH+oKDYuVGzaqV1EotdiIEkFmaazYxhOdII+6HanoLlP
bifilPdvlp40gS6vXl/Jbj0UJQMHiAtSBYQLVb3DbT3PSFhnVuRyRsEjCQEZ2qtreEVeejEmqTSW
Uv3zQDKSNzYoCq8vNTdfLW0DhCBJ048CFetgm0uifHVo6LC3dppCGB2JyddaQO9jlMbxjyGryBu+
gJ4XAlKrA0xlWnCVfcxVxl1BX/pXWCGzCFN5IOkr9MF8uqDjawyeaXpghEhXkLz/Gy0Oy0JsP57N
6omAiNiv43IXmqzEH7RWk8fBPUgzyKpktWKnx00yem4JLhh2yinG/K8vQ4xbFC3iM5ehbjdl88vA
YJcID4dPPBZGrTofZBQW96Tmmp07FiyC/eFtiDSHAAFLXZhZHxER8vkpe91oO9+dm2S8CgtM9aNr
Uc4weri78FLBAKfPLgGv82nF9tLj/NIVSCqkEUwIfhEWZkMmdkYh2HdmiCqAi2WSbBBjEzA7poK+
4cam3MV7ImyI/W4+wXBJppWHVijN0oU2ODEZFW1GH/8DhhQRHA/sNktcEu/sKz0Hr/v6roq/FIPm
4BUCRmQVqQEDUw//jhEqODgRyL9S7tZzyn/h9s2TBBsG9ftoy96/85gXp30TyGOzw4+5/VT+X10e
X2+zpbyFkgiwpPNqS5MkmrGkSPYS7TrH3z6UpNs6EdyF94wV+1wJaeu/Z6EdsUern/12p2jOwnHt
02JcdzC+LLwZV+Y5H6iE2w3B0Thna5vZmUxuNYyzGpcbvZ1LHyEAilXo7/4l4qILaCqIomrIK/e7
qP+43Y0natQ9uIAx/zTBfoNNKZoscOMcJ+ZJhYZF9KiKk/ZKC/dHorTcQHhvzmKTxth4wIGK/CCV
3aP5eiOhFkDBarlTkNgyqxICExlxQ/qHRUcJetpUb54v/Sgtq5gRySAHTeTp6H4o4v8/yR5JLT7J
RpLv8MMqgFrnc9QR6nPw90BBo3UZoo0TLpMCTziE4J3nFwHjBWDgExFgTzgdtdYo9WO4skXpoA47
yQ1SUEKA2aQN/qNfcvudCi2Y0VvNRiiRmzcV1HazFF0eKgmM1Z8YWZk1JlY9lw/BgL822X33xgnG
9Qwc5zLEukUHPcmyyPJgl19ZGQFluQHUSEKAx5yMg76RXi3PHy/qv/nwg1P5xntcqpH/Z/FraxrA
sRTDGR2R3A7WBxDNdnMpSrGfoJDJ6HFmYp195WrsZejdGr/6xzdKNpSYoxh0TNoYu4ehA8Y54SNf
cKLk21qkCIQhCi7eY+anLWvZz4is+EYQNHRx7mlm41kqvOP121rE7HCd+hISDC/JnUKEkckgSQhV
MEVcZVXM8iPCFzqs/AntGESTTX/J288F8vqFe33xMdkDd93F9CrVfnnNv5BsZDJX/j3plYX4xPTv
I9i0nWsLgn0k1Io4ZrN6pEgquig0cfXuJhte4ySiYz7EA0XQf1abK4NBW4IEBbyWO3qjNuYZ3+Pr
O6BeqIpGcGkaPAsBf6JTZBpu11gUcq87OUH0Y/tgK43RSor4ENYlv1tlAQj8vrwtQv7uOgVkB26U
iFb6wNhUfPkvpg2mVrrHNl5TJql83rMpNc/ss/3QCRQxg58XUrTqtfPw4IHYXXBm3X0MWysW3CHb
K7YzG63DyuV4w9iPVc0Q4dvlh4kNWrt1zkPICBOt5ZLwD4BI3/lFkUez8Qzh+3bq4kDCf7T0o87F
GTorUBI4+xoJ8Z93OLGjq3qcN96bouBNAk1nL/jVtaQveWa1y0Ak3/fz5S8BBsQ1TNU5gRp9ygSA
PFdFrEwpBgmKAQgO62jlw/yXyZ9FaPUm8vF+F6T8J2YTLkSTK/8eX+ZDYiBS8AVAOIgbjMgwBJ3Q
Czwz3HUptVPW36RSEmiGrl2qyxvh3XKLmLS/MpOx5UhEKGOvsCFt3Pxi8+ctXlPk2unKkWEqFVEA
ZI62awK0AoNdtRY85k1IFC/Fbmer4j0zwIPKu2ra2tvkr+Az3B9pC1e4vDzR0Bm1Y+xed6xAnDO1
rWiyR4TtjGGysjX5te4sLasIZ1iim9w5qW07CGU9JKbQcEW77Tf61KaVrvDT8NRHlhmzPSfiU1Fq
eaFT25DeOyrEHhoPni+YTCh/Rw6FRpWbH7MjqhlAUT0RynVREHckAyr0BfSYZseYpxmMy3pn83NA
bIdHa3TgTcY7iyv9vGjdkrAoGwjyriPseujlcG75qIA5tPjg/l/piwHExjM4r+QDJLLOhoYJSypw
V24TrmuHZdkW2o+ac/fm6kCfrZqLYR9kJNK2jQdaSI3Fp+LBuJXL/gkhBpWAMm+k0RhaRgcGjaQ8
njARvWt85psyC3DvBxOo5TzHBaCDV5EJxwSmJWsxhmIodXMekOhSQl4DFkwkz0dVdJxCBKOctupR
eXBhivR2FaJCzHNPETPBrO2V9RaIJYA5tRKvlCfOMxdLWvbm5fRlIavd/5ccZeeUxGwMhYNE6qyF
W3jqPJT1tv7iL7On7NosX0A1obfrtkvNBFEYUEfzFK73QywL/2Mj6zoVNiUeVgwO4IfReimSvVCu
M+1RJr9l5hBlwUmdq8WVz24MHaOANbTlutiIRtVBMfLcjl/M1ZZjXmaf/PRnu3kMZ/+DPgii70mS
Aw9FSRHt+8r7cqgZzJ/uQkBl9nNTsexFQK6h5+p8y7x3xuRHr7vo13HXyate00gEobgIM/Ts+Qvq
SnMMxl0CL/x15isz8Y6RkHgcgG/rsEu9Cg3D5N8nXN/wg2UUkzGExv19Ti1KBpVzVwrj16KZFtGV
foTMpnNu+Q9sQVChMdgDREiW3YxtObhyUCFyXfZzQmYS75i9msLJc93+M4mFVdsXuxguMb9nAQwK
ECCipOodyPK0RVvm13MownSaxGcD1PeGg+Ypd1qdaajPXKJwazUWnxM5yDF+cRSGL1iutdWl11ci
8jF3w0CitTu5qaTAWAHXVcmkMDeyxYo6mYIxyF+snzAwID2MgbxT9PDBmsKlCkwbRsIZ6/SkP1hf
ODxmqTS/Jh6t3E+4EJMFXOhEXB62b0zFH+von8whvrXno9PbIMB52tqOxQaLbPYzC5dTE5cztHhw
5eMs5WRWA9H79+mu4vg3QzfYl1cF1h48vUKJO0KHL6N3bRYNGA94nX4dWiceYw2KH+/bf9X7ItPh
G8Hp03GVNRNJfE1gyBr5nDHgieMZ/9LOiQ2n04UbBVXQ61C8HlnPt6WlsxYkmuK3UCgClJVY6cwO
AizRw97BkA3mEEoSGAzDm/dZIz+3zYqF0Bnaaiw2/mg8piktM3hIGxgprspz4HItVVyOuoWBXuQ8
uAtDSOaQi81WLkkK8uCdl4BE/0vd9UzyYamv26eTQhPHH7Zrl4W5GxHyP5odA8h4+jOZsQMKwv8+
mEavltBL5gGCdRmcX5eLwsy1nZrrof4zqZDFJlYATj2KUbxDXlQWCCUlnbNENqFzh7V2Y/LOp4YB
wpVf3fM3x9YwVmvvjJhTUeHuVc2nQoAv/7JriHn7oIMjT5XnfpZdvUyGmUPq1IH/sZ0pNl+7ugT4
GbJS+5jV7DUZtaV25sMrUEdXcGDJCSSRccWuXVhkBEvpwxEJp1tIF2bA9EqWw7mmlRGvlQxhrtx2
9RRceoB9oAF0apJj/vOouCL4ZEJ2NPirnWCdyYpZOQxnqBkr+RxCx7AjmmTQxmI2Rws20ElWS3fs
HbRDUzR+c8f+qJEknQi1on15Ggen7zLrMBEc8qUyYA7tLT6X0bPQckqdd0YFhjwVa7HNUGzDCsVy
ZPMkMlAhypABG/DLA1sjPh63iLjcEM8KXcHRv9/ijr2lsdbYvvMJSsM3bssoQtQfHaE0/f0Zdjmx
Bx7XQ6vKDzwjf5S4ZJikVLRsIg1bg7OcMzsFKEID90BU+dTz/GMnIPJ32e1DabDDIIt1FQA36yz2
xuVaE5AcAKeJYVIpy+iAZNlMu6Su01e8XYob7iSI5lnyE7jThCCg8CavICjEkSrioEaJOSeqZ+hy
4QB/mgDuACeSYBQqcOFGXZ1hnexFJ9XvGXYyh7hkhMEEQNhsltWYCRLYia4e8wiHX5ZcxVjzVUre
JiDSQQ+5+2ktsd7wPHzPebRhNkE6cTZAdlKWQEJyh05ZRM1WZxP78bgob6K+cCkV9ATv2fFehFQN
essosUXqxJqkSAgIMzbjAqXUPctCcf8IYxzh5KZ3ahC21Vw66E03Z8GiPerC+nz1mphn1v7R+80e
ZyfouTptRDQD/kkTP9HE+Kb4p4ApXmY4TmU4MRswFBaQM6V6QolWFxry5qLX0/4m6bsqI8yrexvV
+zYV3nuosi52aMGxySo/w7Ky7+VQaS8RjFdCcoX/eP3HL3QJQOcAebnlrbsEyDhFMMygexM6U5ut
w90SdrJ8n704dNP1vCmap7Uw6fCHZ4DSht9CLTTP7SQ8MQMci4oBa2LOxLCBTLJrqg7pfkfqxyLR
pWoRitFlqFkuAoWBg6XSq1lHV7PKXZDHJeZRAoyiQZ9aRwk6iTMjiESgWYm4si4erDW4y1yngOkG
+ImDa2ZA+4p8JFu2yvd6WXqKZJqIRo8pZrvQqqvztB00xyqrvWE5nB8uOItaVBC4Y/bfYPsqo9zr
YGxszRbKjRBedXi4B3Mgb91aayDTkwHYMzF8V3i+nNLe2Vlysp2XZsPQwJr0Po5VPH2dxJgw031Z
hHfD8R7ZRSeOT6u2g75tgF1j7B2k7q5h3bVu73yaFdobDzilOvArKDiwAIT8sjEgrqZN4geoWrlc
ziXedtiQM6A3JYY+sG0+XKkel8eTbVYuGEMdtitUTKeQ4lXi/NJMv3WBm+MIRkN/RkYLKmzU3Uhg
HX3ogPifX0uCxLvVNc1AaCHsYNjxl62Fsg/ZxdyTfucppOr89EgyNp7XCQ7L7e4KVaaUbijMm28l
tCrnXj9VpLHGjhBcqLgoW1w06+9d2SCRLBbS3TMlAP0BfZSkdGgCDaJ3vuW2fockWjprNID1R0Ut
HeSeoC2kwWjaZWU0JQaugnDQOnLNm/KOAO7wrqy9XhbtEllkcSjoLQnt82WTADVElaVOr2Yu9VdR
oHe0Vtu0X8svta4Yf6/eLu1cIvN8wfMNo8nohLdoNSYkmB/SDPSeqmNyUexxmZhQWgEYveNu9tac
4xdmLICe+SEBFu159LvDEAJgEj6kouQqx09S7FJ0dMCoR7lW5G1i6HTAu7KD3VFcCeVU1StRbwE0
lhtKRxT8xXaKxkqufsa4vikQ2NXUqd85Sn5Qsr/KaHFcm0zyTZxMwhIqNP4DhK8gqKMYVcCQnfZM
x81ulff0Vh3V3HA7AP1jBLY8BaBi5QSVqPQNpHKm2sgpuSZxmqOtWEHyOCQUn+Xi7K4gOpnCJyI6
3T6q6lfcrCD3b6y2gwd6rJyHwwc0chkvQUEjhhGEYsY81fUlcViUkPH13N9dhZOLL8v4mAY946tC
8VgonoQgvhEivJ0Kst7rl0dDNLLl/lRkSAVNXTiVlkwq3NPA9qFIBZmrLpDJDV4f9g7M3YFyR3J3
wQADOK4ghFK2T/QtWzTGI4IvPZ42DGT2DzPTfMN7Lih3G751e34F/YSYkaYrxLO+C+FYo0F9cj8I
pZMSbe4wbiWUi/SXdEFMwMTyzwHGwqCWKHih4HPAAfIbNXboqv4zpXgQ/vTWSmfsD+5FtL+EcJ9B
VDUlg07zRY1agZXmVVXHCCeNAaWxy05aXxZ87WbsJ33JZxLwxanmkqAPBGBsJmWkRLx2zehAzd/R
UAn1gpjbvFKpidYHzU2s6P6dVtETA5t6/8V2JJd81Lw0vyqj++SepUnz0W8eevEiwwk1phvdRY6t
ooHhQNCEL7UYI+AlmOd7ozGJypXY8hdZzFkzfxMC0uGqn7di3oJb2rZjemRyu3dd81MgRkkBiC7j
hhUgahNQUV87LTXv3XkJABG4TzN16nrQZU1mipMEAhpn+0/967gS9mVfO1MXlyIh0k8n9oRyhFOP
PzdcNy6Ui8KAZtep3W7c4p6ZtiSsHAif+2lHhAJnpxJ6iVCah7vnNpXPDeY3fAaz6nMnSM0Vzz1Y
gBDS9TXqibe80Vmu7roaAv08a33vR7SWhElf1HTJSfVTBzv2zDNRtvubBPn7EbxYOiVxcweI255w
qcq8N4NJzG986K6eEljF8hYerwiE8JIB64KreHOQCC2Nlco+6bk/+Pgmf/ERjhUtnL7yFwmhU9WN
XnjJAcyzB7vIVKK2G7vD+rEVDHQSR83SSfUWH9Z6MOXs3yVnBkDm7q2sExXTOR9W/9bYv7g69egP
0DoMGqBFenYjXunzeaWdEWENpcmlU7WgDBSm9qPiP1mgoDaKR/JRed/RBzJjMD44J7doso4IW5/Q
JSARqRMRFLmK0c6W3QUazzUOAihvnBgbYYqmmle74fsvGxHb/6+XnALZ8QBPEz/MkHc8fIdLSPdY
HphIBN2Lpx/FTRrKRrt0inIunC3qovzxMkHxqN3cwxVtNsxSty2OO7OMButiE28dkZa5e5IYBpFs
cIcikeun7HVm384vgORcWBzJEODt4g4Wa8PTk4mkJFtqXd8BiREVvUSdBphKKnY6lZdnflS+ywPt
BfEJt123MF5HnXS+Gvgm7M4rTlAhJ1axFL19wB9PQfy/phUmI+tlKhVV61sGruJiFBB44Zr4A9PD
M5tbZ1mv0Y52Tu5WgJ2NgIArnpipPiuB7jU15yA+EUV/n5wumjfvGUFDH5IMl2oo5Pe/RHGoMgQf
RxslDtDn0dPMZLgy+AQlSphrJ5BITBjde8b8GTO2dG5buhNWL8UakKT97D45KrzL2v/MRQZpLLdu
9OPbsfK2F7vlxPKugs6Ej8rAxVOrQRPixHYknYnrTyDckYrGRaqhclcRutLZf0QSWj9oiMjgMJPf
J1sz9LPSCB1+j8+LgFWRigd5NhRSvnmFNx7P9lym8yLTCVAlCEODZb/hx+OXeX2dc1ADQQ+aID2g
QuH2QPzb+7VfiukcXI6OMyz4rHJ0nRlpeXp/K3STbQtqx6DChC9eN+Kn436LT0XKn6a6SD64boFn
zNq3EgUZ44j0YkwcBt5rc6mL4499ziz0gNUqfuxJ09hyvgApDFtUf2lbhcrILyNZ7wD2C/NDpXeO
kRAGNRDGOjoyBWQEbFleVYw+2z5giBM3l/40HXKIt5Ko/d2MISRH6/pMeBcpUd4UC5ZZk8YlcD5M
dfEJbOe0oWNob4CihLEBSJyjDv20zRw2QENEzGFEC8Rq3JARA/tUfnxODUGnSFdeOYEQGAmxJ+9l
/H5KYjF7elanJllGwMsR88ZhkAdjE5wGsokEKxDjHGwcye/QukoxUTl8RmpBocevQ3/JHTDXRHjz
o/oi26ET7ufFrueVpEbDptHfC75vMHcq51QEsl4bG0y/Q8aPOKyZzsFlA5tJ/rLQhFHCCl6SG8sf
3Un8ebdeju5w+OBy7LqgBhZcaM9QzimqGxm+Ubk8dCfX4h/MAIK7fhKlWVelKEsP8xodbf+lRZ3n
Kkrry63VftNM5u6VvDQVfz5CrWFOUzrc1eCKrkCGfMAwKRGKra2vSlky0OXZD3yyEBVLi47XGfb7
2RGvwDg089IWLJRElsWG2yIA/VMbMY92sWQOnEW98HABAEmAzFj+Ql5Lk+pnZyk8B6NUVQzSOXc8
zLdFgt7FgPOKJIdrb5CB2JGb5VmB8eQGlqTMjiYE7S/0YmpFNA0WcpVbHwmGK7sAWrWfUcPJsPGd
mOY0d++0q4mC3uQicMwVNOIxU3YWEwHjbUvhe+rNA8a1DqzGTznyMGpbTUQ/F9+VfrumaWs8aT9s
W7Q1uxzgaTPi9kPVSCHK+qPJZtDKBA3uTh+Y+Ik/coNFHDCxijmhZUHfMKPN+wmewIOFQP4e5QNn
d4tTM/zegh52kAoNILtwXoksy7RLBFWo0/hvKdTE8ePBU5SiGDx4Lkks6+/HtOVxz8bJ5/AMjqjT
K03nkG3iUnlXG3gRvEpgVKX6/S9/tRuxdVk0k3xjTeTzC5KbY68MbcWbGmizd56hv8Y3pFBzikV6
crMHg0C+Jgth7i35KNLo8I8YbOTE/5FJJArbVzuPx/k+Xy/hHA3uOxYdfbshKF0Pav29exERTfE1
6/pgtCnfQc4PFqoZCJApbIHk4RPb1iceku10cYWifHXXGsbr1dLXzO+q3hUd0DQ06nqfJN4whrfU
CHLL8EwXaKj0buNerEOXxmzNBi1INRXFI1RYKhcpMvt0SQFyUtVDgAHWnQKCxNygdBHJHrYC5f5U
xmoW+CArkUxUsPb6TN0kP/65PbEfXXumrb+cLZTu1fO0mXj/T+BDRyV+4cPmRaPNrIydJtJlxoCH
kuYMJi9SQCos9KJGxRwqUnszbc5+Zn1jASVGkZjntUYS2tHe/DuIrp3pqLGOd+THs31Y+0C6V5WL
pq5ivFqRHUC2Au9eIMVvjo7CWDU2TtHIKM0+es4HoYOLSTPDoqqCF3zjie6mfsyJ9S5xZ59QREP9
rsBHWrwP1VqdkmRnnDdmXuKkxX1rEYWVrXyaYoLDooRfiT3awW5S1uBvMQlvGNOw48bUKuGolsf6
sS96CcS7kXTbjOVnHCnxUvfFUO7x+nqeHRZCUqLxlL2ugYvaWNWl0SPf+bpotcAROtveEQhLMoKO
eIqedk8D4DLU1mOtDVTX9IGMsXW+6P9VEk6/rB7WdwoRaquuMU5KORDOLt0cOGdKH4GPnxgv+/ug
ph2ibtDzZASmI3KtJ6z1bfw1EyPQkn8iLG85JbOOKtko731suznzH+wKpKU0c1I1K01jUPIwSl/E
iz/nuCxjFjuq0pMqBNc8ckzXkQ1sxZDRhe/FhZiNtC5Q2ndYM6YFz3D3OP2+H4DN17s2sZoELLQE
MN6plhZD6vcQDei8W/S5yKdQsKuXh+HxrogQDYaOGUBJ2S7bXpYgyOqBTN40VA+ZfggEX9BLP6ET
3bnMPZiKz8RBggH/i31cFX0D9bU/7crH/7VRzvDLqdiIMpRByU8rNOXZS9jdo85DXJSsgfQiiySp
XSktt/ZZZ60eMOJGhfo/WyKFnFT3i1UFg9/W3ylhMMwhNQFFEdC72pCQiTcpVRuswiOEzQASuTGy
oNT3nV69q60DfQo1osUqAotb2y1VNFy9PYwy+owRz1jIYccsqiR+hS7uBl28IJcFWlQdwhxg9VAC
PyrO5MErxt740dJ/m3fYc+4r2/b0OBoOLx4iOVcpQ84BqaiUYqJnW+/Sqc3c47dgTVSDZ1HxBSjR
sSaCry0kEoEy0uURO8NQwiL+wSm/VAthWDBScxWSunnK82mP8fCyLbIWQv6Gv7bc0dQ2Ie5xTIzF
Hjr5oNCXm7zozHTl9JATirwd15raopS/M0JG/Qko6n+oyVA/hQhWb64R5xdX+h/Pgckuubxg+Ig4
lBHY8FYeyx5tN5pG9jvVt985WegHAZ5UMM2hvESgB0FVFNedmxTDvzD1/XtZBUZTRasfPNjcBTx+
cIGeercSzDkgVp2q457qXdexPqlOoHxTvOHxFIZHUwt+kE8lj2eafUxIn4MKidJP6K7KWRs4SxBU
3p+dCRbecm3ukFpKm3MA0IWRYSLbKKJKcvtaHSTqpYhYEPlPckU2W5+K+TP16HDcsqg5PjDrrZXx
H7a0fDziLBiM7jdqgnNUMSZx4sAygsfbnJ2uHABNGSg10OGUTYrnu/kKuJXmyZVRJ+WieSHoDAy7
78WABOyZiz1jIbv8GibQx1E2UA1GuArNZVHdzwBUz0TyTTZbbvKX7iRR2hTlsTzVynUJvY8iZiOP
i4xxBOjkCVjiYUcDSuysUvbF/Va9rsE8p3Z4P/fQbQBLoCRS/e4V0aU9KhUhhaEsWcPGNsfU2Du/
9nWG8R5NWT0URzyxBahwN+Ibe9rPZE0ZMKYSrn8cdlLE+OWfTI5DWcW+yhpCcy/MLLamN0hnt2xP
EdN6CvoBj+9sttc/Fc3dszM3k2/R5jvB44RU9JSutGryWzcia9tLUEUGBUXLyK3ilr1p8pB62sQA
IotsU9gHvLEyANXFmmiPagQSD0bcyJTNc5NAKcB22Q3vXoQMfkL2se3lDbgXukMgJlRo4wA9jfK8
hkD/QMXKtvZDv4vKS1p/6I5Lh8Pq+yRhtPrYupZukHwuGDeTCTUp5LPdprRdW0GeaXjZRh4Ac/Kk
1laYVgU17RjKRjBA93hJE9xPd+fVr3sIDw88FZ/hIV22ID7NvP7iSCWLs3TjAGNLLu1bQ6NJAg+s
12nvQMPwSxkoruc+6o4E8z6fU1YrfypNbkmp221GDveo3ELs8871W0ALiyyYUhSgqA7qJWrWucSb
xnNGp2ujO2RbmOmdxN+WgFtayncNoi/TipSMqyJeenn4SPwElmgK05icWO75jGq0y9N336uuYxIr
UrsCqVFEXD/fk8yUerBY80kba1yUyLzYYHN7oB6zGrtIsKxwU8J2vluHGWC/zsW+hRLOHarrbNe0
LrjM50WDhSGM34V5pReIrzLlD8wMo/zCfuwuiWJmHwdAcukhXBNvHAkdUqzcgceBR8V6hA2CQNyl
uwV7QlQl4WulIh61kzitMLAsqn4GeIL1juU9OEPZOvKpnz6/H6i49uHYaGfU9IOQ9pjAAPcZnnB8
xACCxmdIV2r69r9ZETEffNT4JGnezNtL4X4O2IYJrjGieSSIxEHBIjvEMERB3LVrQoVKuViRnnR/
W6jZQHw3Auc7bjaVmUL5Sg2Dqu64j5tUbJNz9/mliKVPgXMSV+h+a0CNaUaRhryEhAp9yc9hxDyP
RRkE/zOOp92a0NsdBTjRlpvJExbLkZUCPlibgKqI3poUtT9GDNEofe8/sD79kjCwrZ0xZvgJKMh9
0CUnVoQN4GbGxzybTXnGldyF+7BYwlltzbK1gnQ9mdefBMx2EICXGIDqh4R6ToI6Ro/IqCOI/Pek
UXJu/5yTx4Q/nZqVB6OMqQu0pMFosSdHq3TXW4h6WVXAr0kRJDTSPnnpDP9/KHbF8etyK+KPc9mc
vuiU51pR1YhTg9hVV9+dat7KY2q8h2T7RU9ql/X5Z2S3U643ACzcFcsTGRIV3MdMXzL/a3k3/lWI
IUcXJ9xc+ZPSQQRjwFpgks/d9tvJd6K0eZrmVvDkggCDnDVnMpfbzUOb7jpUZJeLswHMRA4Li/JX
opVZj/PGsUGTsZHuDdGB6I8C2XRbK90Dl6wZ/pkZdMR0NKddokt2G4DMNo+Y+VwgpZuzBkaMTEnu
t/YtmFfXhuZr6LOKYGUPVPSPlFvUUV74yR9S3p+QXHf9y+tcmaWzu9yUa3vkxaWbBfUVXIA91X0t
3HCQUrQRtjMomnTcCW3GYWTbTBOSZR0UjrU7zc5R1e7FBOOIqcWn93nzdk4N+O+63KVaZTWciJos
+9/ikbopbAmYgjq7Eahurs7E7I4kRaZO3P2A7YjttxnTK4YgC71aIHtDDwWx+9KAg785h9iYDjS2
YxA0J0zd4h7myrbie7QXt6XH2KzwMle3DmdkMd7hjgcfm4AVJOObZXP4GWHtQmGyQbGK/HxftC/5
kESGXMubHu305e21CuTG5oyPHQ5db2+Tsjpmj2h0mXYUK/t1gkdAw0Z1w8dnQCcEBxInAuZvUUtt
x8DXTbBlzCrtM932aSCJuMx4rCbNPh/dn/UAULaPLcSCxHk6D0SXP843b5UYaGNqrZWfPPR49UFk
BoIxPXWCoC1LILPDPxdSbZJvWf3F60RMVfSH8GylPoq8v0x9x38K/xbQzzDzGb9Mh3Mqr83Zs//K
fbECxhZ4xZ7ZU5p9UFCifIxbglw5xNKp13xsMStpE7aiH6KRiF9BBgckdqhX+yFW9HTYKqFsk3z4
fAqn/ycIXaFf7srxZeH7Th2klra9UMWdolfVeXC/hJGMNvAarU/PMGu1R7QC1gUW7G6DeVh8c6b7
NZ8nPcH3JxnPB1gUwjGbAmpNG58QmqEHVvaIkzGKzamXdsMvDGv5QuFxcFDDThI7d+d3knLyGgNL
9aytedtpr+JKCD6g2HsXJNCdbFDihuxO2oGpiUEJujrH59n9bDeUtXBZUaWtfFaDdIicZFsJ3HIq
7MtT/YtigkJJvN5Eyjg2gZ1/17MtKg14Riqemvj0iIKcut8bHspN3WV73CPw1/z3EF2PDMdA5PY+
bj/apY41dGhUkXolUKVLA33FecnbH1ippgJZsT4fzvF4xb5rmsHjS6GlYIsQNiIkP+788vhmGQJu
+ky4OyWBaIa+/fGaYLcqbjG1bcxnh1Hvn2dlSEogF1fK1vNVf+e7zeoAFhqAsl7NBwualosPxikj
qmsfQ7tN4NzPraPQs1saBgWS7cUgyRlo5OhAo/p7sdzku8HOyNiDIh1s8UiBqtC0MdWwI4AXIz6v
y/ABE5L8fe6y6xQaCOp4er8l6v+vnQWRlUN3ryNv5hpnnEpSwmKmer9aCz+UEAaNbITsAbK0abm/
uMlbrvO4LF2PkEZ3Y/dEUv1d9/Y0QeYOXe9ViXkKbedsBBWXf8erUIaLvVZ9/k7h1/2va49EpKlX
3N865elx/0Vn9IvO0sXROboDgXrHjzSSCmAjoIMtGkoNRyhuAcnHhSuGHpHqqlsn+QRJFgFy5Ubl
VNx6i0a9CDHwQ7heajEIjwpQ5O3rh0eU5DrkcUHisaOu08za8CU3Jd+B6dRXfolUkvaZti64pfX2
Qs5NqX0nbGSo8B0qpbiTzjXpdcFZ8gTvHBknAn9BYX84eAcyjG8mbFqnogWkcLG7eZTe7rpAPXYi
KOCb/k7q97LrV9XF+nKPb87kKm/fOyNqhjXHu3xKzULRtD1WX1JqLcQD7xQ9eMK4ncE0UdIsiHi3
Go9EQMdLJB2r0KoiRntllCnzoerHXfwUfqyl4a15TUP/jLLgH+9VWNiv84DbaNfKfjtLHLU8HRog
3nmrMCMcxk3a7+ns0OClxzv2nA69rX3nTZENexQWRK5kH5096Zo1OT4jy53Nux0PGCDlm1UR/WG7
bHhTXePYreS+0mdtE0nsGOysutmmb8wafIo7cD+1qwmadJ1Ohyeldg2Mr+0g8ot+c0713iIMAZA9
Uym+UsT+ki0q3O/KLhlBB98zLMvR61jbm8m8YHjuCLaj7xgPdU/krtE11+tUgRI+1Bv3uAa8d/W9
07K0vnMYMtvwBkK/kWnzkMjyRwiHuGAdp45Mg+27MYJcy2sW8uNB9XepnzbfDln2l172ElgjmhCC
aIZmPm0VKr0QubqXFuooEiseVDJ7j9qXxlGvvr3kxBj66GqFIT6ua59fbOgx4mX9LffAhEpRBwLU
4pNNIR2CAe+nuobax9e/nV8x+tupA2bwdHRO6JoXjUld6620qbzv4/fbt/PqL2zd2Z+I8eSQdojw
SxFCNEhJGv4IfIfJfCic4gWuUdBkJjN0W4C6a0d7BikdeQonqZH98MlKdGG7X8aT//aG0D/OeB4y
PCbr2VTflOdjr+MtXAwnFgz0tmVYcCxRAp7EdXkLxayFEfzMv2bTV0Y0WcGpMxxU2qGa70DX74LS
30QaM4VzWXL+omTHIjgConxW6UZSDsdmBjIosYh2XzSthKmN0xgWzTt6/jEO4NeE69+2cpjQoSzZ
snOABOrAySNKiuJiN7azw7h01Fr8SVbNFsEW83+v7My8u8gINHaayuUop8+zedMfuLNko5fvbGKz
bKkBN+mCVZj4Hj7Tct6SOGkkH6dh37dKVYgI0wrKT0R0shYBE5C27fh8KDvr9hTGW3vQhBqwBeko
j5bveZsZUXqiiu2CSSb/UZlQG4osmG9zoj4XqRIILXyMd3rAwS+ENuD/Y7f55ZuP8T9lXe9QOd96
1cDBd6kqv1R6AG8FPb1VxnqylltCF/lVdAcOsLc+J8bYxqqwQzIL3XJGTxtbQXb7mw0y1B/yVcJa
VLmyxiMO0poBqvl72T4bv9wijINj0SHDGUH3h6rJjgugsz0ZVQiu6xw+znlRdVzGnVrM7Ks2LeKY
oqkogcY4YQBhoVpxooLZ9efbIR8yM2XvBO6cqmBuFebY4ON5DryXhjaFRtEpERTpvpM7A9Nob00S
7Vd2/oVe2A6TEejpxbbyzyUTnixsbG2ufG3m+a1rwKM3IMsu7x7o9OtmihJ6QtKJgvz9CfBYKNNR
+voVfm6KqHloNU0J5NY8yTfAG1HDlDFVSIloTi1V0JOnZM3R5tz7iy7IjRK0uPuE/UFjqIKS2pK+
b/YlsxgtkqJV4fx41gtNEusxlPmFjEPRkBO+n5MzPCJ4ppVK/R2BXCYsq6vuxQpacSAbIF7uLwSW
QhE6UYPmek0sENymOrjwgZcwZFVy2Qd1T6rTk2rB/bbBTuE9lkr6apuxBemusBI8GzMsQQABPUgy
mxPAOHISr2P8E/abj/4HjpiAxJBUyMQXtmy0ZChuz7TsazK40gBCJNj6QhkSkKsqJlrbjrxoQKUt
nH8DIVCCavqEskJSiJnXVis2x50Bf+koIRt1P0VY43sQ2Er4NqPLH3mb0gC6EJRkAOhBS/67+kYX
oC6YFk81X0BtZGx9LkgVaTKDC+aozC4AWPUT6mzFCxEaOz2jdq1qaFcy82RQx5jyON+9rP7h2FpH
J4QQwuOq9EtTnM/6wgk82QYx1l45Gj3guKtfTTYJQYCn+Eq+BJOtHzM5zZAwL+B4oLKr+pdY6/7m
9qyFs0v1Ym7Pgt9KSrjBvyhts+/oyo+BiTMGWB7fUYmA3/1gPL6UxKxfkV5SOtpzKzT+WYzJahqq
xGnonFRInM7B/99yVg1x7vpeffki7RMDAFpgXHNz8JBYSGCQfLogpDJCCS54a4FdBnZPpW7a+Qet
Nj2u4jMh/jr24tJQnk969zyL1lowF6XYrFi83G0UMO0OFYskhljIJIHmivysYjVONbINT1FFTgOg
tFs7Jc6R1PBjmP79GQvb34lUITbFQuiOBrxUYfU0sO4yuJ+5KSqdcOQnccDfCIRqoR0f7fal72J0
k5MifmFJJB9L/hl676+uznBJ8UvktJjoFbWIylf4FpxjyjggIIw5j6E0uAn6vUXYAOm4EenfGi7b
U0EoaAzdRQQKQC3YKE1uUuVofv7JyRGt/QaFj/41CV+9pW1a1SsLH27o8Xrb557Qkc83yuf8t3rR
fLNf4FpBZQEW83lSQBefd1GkG4c4hKzq/3d92ixv6wjZgHwQpOuxU7UK7x1IZdVGRONNt1EJqsyh
S7vRmF+tfeGgvaAhk4NiDMALsd+ZzZNCDAZlNpfsqBSN8Vmi2B0v5/WiaFFfAOspqG/mCXLBODxH
gPZ2HFXbGtLdkC9Ij20V7J9n5f1E5i1PgUcDG9TieGVQsrP3lywjk9a2HM2zj4c1HIdcf1nM7D0p
ZR2lb6efeTh7I3AeVtN5QgC4oNfYb67T/fjlHM2hF44omZUHY/yXcOhq80Bm1EgC/BPQLFuspqhC
4x5RGwNOE1GMTVHgtRn224OODEBYYALlLvuQxlRDUJsQVBPTVEMrFxAsG1h6uyudGtl82Signn9G
O8ygLS5YwkRkhLg0oJtvZZbcB8LUMZ3uPSm4Fje11neBaiiUio9mcmkOCB2P5TmukoK2uZzxJrmU
Rh6sXNangOptFNUBn1K9+Xbb0jr8xeO2RV00mGlusIo4ZmzfgCP6Mi9o/XU6rfjZGG9FoRrZyKHX
wWRTJEO/Nf7wKTBlwX0nQoOaPOxDa6+Y9CoOb1h+Qln/8dqsfcDplXKv5iQgP1GzMWHwKL2d5/Lx
SI/pBuGsYVigrBqH5jVahnTLlZ9Q9OGJ40XhcjPvbKbsUKciQs0JZvUEkrnua9FOyjdJCnPxsGAt
KbWCzUjezFodjrE23WZgSSoYkmYxPXRzbW2cEjNaDLp8UCu+1dI4l/xiYX89gzW0JzHpfc0EHagG
rJnFeQiUP3om20q1jHlNwFYaUmq8DVnPiVOKmnnK4nyuisflCYfQ7Ofm48HYBMkuJg9b/7N4Xjpm
DQo0R6zM0R0gbYNxodUnL2P6v5xu2z50KzixMvTzE7Mn0XSDOsdq+Tf5OK2D75YQ1TZtYD/LsXeV
vf1iA4jptayMavyQl26sj2hK00ASC3AO97CLztznc8/QE/yzXvE6ZLkC+v8a3xmwurmX6Fda+W2o
qws1Ap3XMI07dm+mVTiDlpyauJ4NQC7gO3qu++utVdzfJfDDpPsauI9OCefkuJMgx9PD9eSjc6GH
MIRytPnBXWLs3NSVHHgA6+FvCnBn45X/0SoCtDyIU4xS9UKeKg+kSiMMyMEeVAbDvkRpQZSIE4Xj
+ZbaR8zhEUpc6r0rKjjsECFLuzCFRamPpZoEIAF2kIXHBh0oFLyDA9JbLS3QZL8QVusGt0GilA4f
pddK8PYPpVSiMaK660G8yH5pnaeWNES1cJwvmk+yLUOrbBkdHUY8OtGX4OfifZ1Z8ueZb6EL7dz5
xP+QOJumZudTQN0iT9XnmcZP3JYzV9MeAZQbzK7NuKCf5RReJBx5qFR31emRwBhsXdiv4xko32vi
Uw6eEnPvudaQf29mkVT+dAuzS+e51NNNTr3LRQiH0RelW5MoEP5qXvXoDnXVKJsFJ5RUvhz8izPd
GdbHi2LogcUsL+DGKPvUqJJvMOi1Kec3rBG0abmbj65Nqo6LC8fEzKHYvI43x/lTDR8hyHGVnfMW
6uTCpCZRY0GYUMwil9sEJYwh2bU3l+sUlmiOxHqGtRnbtAlrxXpun2vs1dblNee+lOkoLTKDZqYi
zOa4shNobJjLfl8NSqE/i3pxp5e38RpdrFRVJoo3ZDcGeoq19kuUbOURWCGhbLnKEtTCWfhI70Yt
JCIsM55Jaw1l7Vl6E8cM7k9s78NFy9cLCMtns+7Ky3TEGJ2+OrNkKknttCRfmszEKS6NGPPuKNSW
uVPsZfObLbRFtrSg0a+EeVouidp31kiTleLtfEF5G8AZgso49jI9sE/lqziYWYPHuMZmK88d2sSg
AUTCJqHx0UoMyBtLDDH6k67ISqsTVcMfqWr3kWJwIgjA3/KlBngXTORQUGROPT/5GCgF1MIB/UsL
wIBOZUfQQHcvpSRFtKHjR6wnF9rtqpepHP84MvZjZHM82/5QX1ZOwdilD3Z70TRQVI3SoSGepJn0
4/FyuuM8NSLogDeDss+Gj2GIiSeOlOmaiWRow5SI2NVSGIcj/K6yD1uJozxpTfM7RDM4MnXV2r17
4S56+JmqW4tNwHGYckiVMNioAAXhrYYHcFrsSv5+WDwEjiG6KpqaQ513dcftwEhOKbni5CbVsyPw
CHuDfVO/OBeJwkiaVY6Fw4AFGuXzqd70usBzdftm+W+XEQEN5F42nzOZkAdvhZfTJmEOtrtvdJQ0
uXPKdvDb9mZV8pve+0xeEmECrwZxW7IIpPmRk8dxx9ExJ5xElquYAw634PxZCUQBpsHEWiGesAH9
DgeyefHsI45Qc50x1gQhs4lfhwbQqOZWeixvBH4mUAUO9hQtn/8RZl9loQIVe0A/9fvrfxUkul8n
uHb7s12OpJyRvKs6pEBVDEluOJoLzsdI5X4ftTEwnAtZGXHxDrgSAMGuvlbQZGKBGeGpOMx8f7eJ
VBt2vrDK9qHc3YrdDd3G/aexh0GEhhfjPq0dEfde8vvei+Dd+8nz/lhZcVi3UKBgq2dbFhn++bUW
Pq2ED721uSViMXhVX50ZIrE8tPwIhkx8318ReVgWi35l8G0MnZ7CoVq9ovArLAu1iylrnmtmu3yc
LL99/K9dXGEnlHFPT9xi0zfjF6X1bYLWLNoHzHf65R3LhZwgqd1yu8+JosRdwSjfbSJx7EZDWrEW
quQgtXcItHXO0j3bRsMMcqaSlnFkCk2hjcoRSyZV5aIIH4DWz0u0L41FlbYNLoIXESByUs6vr7LV
QuswCYxWsptwMQqapURhbFz2EJj5OmuwSH6eA2B+Y2iNUD/84sQutIQ+LXhTeYWvScpuouQTgWNG
aomKUNkuG/S+lQ90636GCQaMBnTf4PWboqlHVfxDs0pV6NRbvy/w7bfRGwyhgG1LMtcLMOA7c8DV
QKDnihn1Zw7oOz5JfaUfbcEDNydrYH02RILYlSkWh0SuZayIuiABq9cKeqzkF5drOWam3orcU2mZ
qEFPpLfx6xDVY1rAYK7LXDEWsorYydeAwOg6Q9e/yg6mDqYOi+CozL88Y2gXFPp6Kn8TjMMg5P2m
upqtTWov/0SorJQtg7VmAcCA6maG4LSSF5OYIO+mitlbHDWkkHycWMQrO6JP2Fh8HStw1Yafjz3h
0p3inm62n/SzRMRxdSsVOhfcQ+QOjjmjZVbZM3FLTRutZbwBStiOwoX2wDego7fbIjzwcF/4bEPV
hdGkw76YvRnegtqu8qttvmpp36RHncOXzOxJMRs9RzORsdoQokJLRLOOlStLZ5tLI0LLKd+pWPaO
gwZsR3ZjkvLZ/vigSaYTP3Oskco4r+9QQfgdtiVwc3vrltxs3XVFd4HbSZSV7xo3j3jsAQdcEfzm
eG9/4iF773yZycVv+z0/vXgp2Rm9/xJVGoYWCd6lYBvHFTVVqgn9XrN/NsOYNn170VpItebuZnpc
uCyj25uBioi6HavZcKGYYOqZQJ6ZEI/MWtVYYgC7lW7S9j+uwZimCquGARXxlrDN34OGqSBvRXzZ
rG7gURYHFtG4zzcg49SS8TynA275UEJLioG1EbmEA44jP3JShw09IAsOB1DqrDyDLMs+MpvhBNkB
KGexk7LqKQErfSZFpHeF1rMVvvKFf2S+HeCA/oCsDTUTgk3sP2z/0KeQ5Kig6OtEQfUEG5ab7gyj
Cqn24bDfpgnh234CF7kx8RQPGdOT+7HXIeLxV13GiolbeFS5L6XOTMhTdZlb72FihV815Jjf2KSq
bQVWDde0BRM8iF9o3EHiMtKUsx2lDwZBbXLETgRAMwcWN2RjM8CE3APNYXOzsa6R1hmGpFO7ZRAk
v6pG5LhbQ5FPuIAYAN/NFWKWQVCj2nzeMbTaaQfqvv37ahXvKGZ7MvW75YdC9rDHzoxdNmOMB7E5
HVqKA29ws6lA5dXQhyVjjwEV5PVvIyJ5Q+/8u1YAMU7bfmTkQhEcY02bX3+9Enjn57vTfmyVKPby
ggT8qTFfTt2+i8wNbM4aOCGBzXnd3rxMVC+yPFhmDeDIFzaIKmnfnbd6awsZ08CUZ8bhakmm8PAG
q6xGRLE0Wxf5HaB8bDw/NQsgdFYXqavnC2QVmNb/51isXYn8Ii+Su1XlUKaNr7Iz8mgt4W+MuRfW
VMQ9MUErVlo2CHG8T1SjikHVOiqRfpI8QId3fkat7p7Fotf4XOMvsz66gRshhzosmp0ECF4Tfn6G
7OVc4ZfXq9ps+Qu0zD394mFE03JqKa/hQKLenBc04y9Wv/EpgqK5csCtUoFRe5h16wKF08rxObw9
soU1Z2ZomEJ08iKTvR+uPJlPEV6c9Q5NDSpdhkM0KZYudLu31MGjJhSx55AVMC0l1tmX4YPQfA0Z
M8ok7Rt9PI6swi24wb3/tA/EX8bMSpQ+QYsy6uegJ1W14CTABYOaf++gwu9xKkgIM9vitJb0Blox
r5VDk0zE+QANDi+5159U8BObAi9mRnwd550omibXVWRqd9dIEHl8gtKztNKq/8oqYMr0xyT6HeGa
vRdxBjcSum90WyPfVgCZL63xtUCdoIO4WVn00CTziBUXz5gdyC2kmUXYNQRbE53+cb1OV88kQT1r
0k+iJDedBKLQIG3BuXg4MbHxWCOpddkF5VUw699+02bih1uaOzvl7O4X1cn12Y6yp+dnqU/0yGIh
Dxo5Xc0QIgzJUSJ6d+vfoKwElpk6pCvXFEVN0QNexpsONh4a9PKUOPOGr5cpivX3Y8eL2Jl+y724
K0liyF9OZpMNvYpk36ChRbQyYIg2yFOCu86vTLijrgaYu8fNexCoqB2tsDzBK6/NXS7jG0luRtjh
+3q+k9UhS1puuvtcyJ5gRUxckSAOk+PvGgAWOdhBeDnwO984ffA1pdJVpNQbwaaaDGz+lEVxXYTJ
wCkUX9TOKhqbohYJTGRXBrjQQ9LV6dKDqCaeDMCBTnwlTaEWSMCTj2Ma53YkgL129Is3VM0MXTH5
Zv8ul+Khn7yD8uv1hpM1pWNqtJmOeBx8Pxw43Hal6EeooZljlTQVry9RtQ9dDtGzKu5JL5w4wVSg
HHvOG+fHq3aG5LwM0WKPl58ORPFwMTKkQqMipWdgg+4TbFUbWNDfIy1wnaBA/fwI41vu9ximoPd9
q8C16dGtGFuTGXHSIpvQYNY1LcBfWieBwh5r1IlW1hVz+3fisxR8goO8DiKWDIvvqIGyPLIqRS1P
qoqvCCO8ZPhUgG45wDbEKlxLSgi5uX7K2Ip3oFSPMNMucj4QGncVaarfGf6QlTCEK+cP59nBpFhP
7Q4QtqpBGGoNYU5fzyc972RJDo66Yl6t5SWw09snFIYHv5FA1boZzytnRTGylLdLHCQLV44ejbbD
awvAi+jq39/H1vSdRquhkGiJO6NtgDIF7+Uw4rfZSOyY8yC1Q3Px5tGHMkS9L/N2YMQrdUToFXEg
HzBXs4lRWxh9ExzP9bDWzqq5DzmNY/ADQSqYrrThhjzN/2lvX43Q0uj/AmqDGpI3xEBHr1ynwWax
UX6Ff1Lo9uxK0HGBWb9Nucj3mz42RS5AFzU3ti8cZiJD87MHw/3mIV7n7Ds/WK7wU707GrHkIcyl
FjWdVdn0lVl/Oz/ZUCiIEhXkrnEt7fku+RW2VXq/1ppqTh+iS/e709h+OEY5YlJEYhtetpVPdwhw
7P+bKNyTy+PE2h3PQJm4Gj3Ytp6LNVPmPyH1ALlgOdAUs1zjXmK1ZvIwviRbPAw2Gz+o3wwN9Yba
lfs87CQdt2pa7rBYhMbBSPGmOONFAJrvqTF00DtJWqDXXXpTOu/LYW90mzmNp8nenM9OBrRyoMiC
9wKIsFVR0OQT9j3NKYanaYp94N1T2fbLHP1fHAjirV8DachM+YmIPGktkHMRUqb1zEcsBmp7XfU9
+rTJCG+IIWXyfBCwf3GEAAdTKLUhFbOJMjVWtxH/XV8BDojqdgYVko+0nGzzp+Ifi61ujlN1Qm8w
Ud7RGYGFEBOgGa+Kib7WVjGR+q2BdCUd5q8bgaLKQYo9EY+cYEbOo4WpfJRw8Ui3Ntz/9DUENjFe
zC8osc+p6rkyB2nK7+duYkAzUnPz3BAFu8uMrrxBpzC+28Utchbx1R/9qZc6NKdavL1KsrgLKMji
05zjgwDYX5n4bSVeL0kNEIkLg9egbpgum54E2d/jWFiuGKdWgG+FG8mNmotY/HRdKF6q/p6YKriG
Ly4sfutr3KuaWzmwxJbeZFpMfSIMc3WJf7jOHnW71/8/lwvzlPOFhME5tEfLSTivDVrvOobWPhPJ
M5gseSrPd9ozJ4fvI8oK4IIrrqpdVpxJsP2SsJDzFDqI06x9quNChpCmsiFbwrNlmPNtaKnMNZo3
jJIZZuR3NF/zyUQPNCw9kk07qYjPW62GJVx6nAgqbbKYNDXBl9h4VomAfIrtbg+eupXzXrTKZ5Ki
VgWP6lFTQPi4xrLg7UtLOW7PkyjEzasj6mpHjTZqsB3wgvvbYO1vzVsy1U6wcnPF7L3WtZz3hrSV
cNDjMMhM0yhLWDkVwFNr9sh/oV/wUP3An1ehR9X/68PLEVTdOfaSPUi8OlXX8v9Z3iJXowKTual4
RsdSdciEPfvt4yYyHwPr9LcVK+Wm8igx92NmTFX2CUKhYWeOk2dkp6fHS6rMeqRsLoIqH5hN1589
UUVaaRUZp8lqmMMLC18UkcJyGZNW6B/ByVQSuiVHwgnDeN5PGA1AGEYNueDwKa34xzZvhzgoHyYO
si8rlzNbcttyyGRK7uEstfnjvtXDoj+yID8C5kWV40z19bTb2LXjw5TTs5B5esAaxghblnEJcGDb
E8DY0BKMcPWFQEKrk9qHLaZ8wBvDFGEtVI9lBDgEVqjawIxOjV3mMqdjptps0JvtqpjpJX6yivr2
EYlKiTMDulqgjwvtjElZaBva6E/6BZbCWqlzDTEevyY9I9qLveVFfM0gcKyVEshblEjIIVEau+/2
f1itRRN750BZCWKs/s9E4qOPbrYz7KE67w3FGnl32VM9/xhyjftrJwUqb6UVztyc/az/lCWJUUgj
b4VzmnJFaS4i+8argFFNAFAbx2k0TseEjhXkS7rxMuS2PGOh7jKMgn2gQzVdRKlZDdAyGqVSYWto
PSgmmbXtk5pbnhKkwBHPac24JaIuFE6MpUZ1CgtWE2gepa7SCjyXRLVDRk9Eo3/X+2Uhu5swrUo5
MNqMXEMMoptvWjlrenEmsLQ+xEvMgiVijSKCUc4ba+xSIpaEePY9K1lvw3Gq9JT/C15XxBomRq6t
30PRSWzBce02O2jW6j6W6d435/Zz3auGML+KiPZ4V6azNsFQ0UUGW+hrpP7opWQysOJ0DJhSB5di
6cQybJxMrN3BtMQ8vyxoRRfTxgqo9AJf5v7Rnt5uMNVzMoxiJo6dpe3N0/vw63zPpC9HSa7pHZV2
HmnwaLu/wKYkp+ZiPSiDwipt0xa03a6OwdNCWBLbQ2Kk4EIIWoZ0P/jDh8s0lvkI5R1+C3ulh8l8
M78DtYCs7mMSEhUGTqRMrajwjrptrLg3O1IwHxYHjKObbvyL2FUbJE57V2RjYQaOGYbYPX9Ylm6m
f+kjIUEgAat+clUE0Qeu5AQUrS0nmBSBcizW9Rp24pjaxL3rK21LYpJvuVpGLqfC7mlQHUBcFAbj
i1Toq1AsaCtEfeN1ZKygYkUBblQVSBiY4uacBrD+xxBWS49QwLML/6B6ztOC3jmQ2lMjLYlbFahU
RXySBWQ8trsL2JllT1W/LND55Sa1KNwn36IxDGekJg8t5sGkikDJINSp/NyiByV+p2txMmrlUSlt
dFPWm2LdRckBjqaA49i13jPypFrx3z51xiquN084oJdu7hw5dKS7EE1LAxCkxLB0VlW27RWDd4xP
J41IHMbhaE0n/bsIHVeTOPc1DBxZF8ULds9QDiP8TlsXCLl2CrWCDAXBi8KROzyNYS2NybQsWbID
vWbSpTvl6Mzgpuh8w5HNdKQIo1e6G5pHmHqRDOLcXhws301U1mS1aK/yy/qtcG+1B706o9f62UVf
qdo8n2/8+UGcA2RrHsy01r/P/6Urua2MXXF/kX6c2jYr24MGImSl27LTFuWecX7KPTer6jIVUIW5
VyJExm9HAeV9UFJNVa7jvQZnSyrT3jBtiV/2ex5QnxhTLx+kadhTCZB6+Ls/BN9MFagMHypMrzv0
++MeV6POg6SGildvaIXmm5lEYxRGh7h6JUkJgd2rfk9FcwhPf4qsaaJSyPPiLLOxuWcXGu0GDh+n
lskMQFg4o+gya/eCQVzXC4FLFMM9um0quMcpve8+sorlba1pAcMd2nxYTA8WC/UE/Mq3hQnvSQOq
qUo1y/xbz8nPrb+LdAIz+49jenYNsVSb+uhC5en4NtgA+my5lBy6iIq4y6NqMx5USIXc59UcrBkc
ESyVIzrC+nBjoxXk6jIgxn4jpkJY+2/t75jhTBcJttx+WvtqR5Gj5bMb8G2Bvzqj6Np1k0v8Wv4I
QYhhXsJ8Rq48s4DPtEtVGQ1qJyDYQXpbC1ayRmi4CZhPBB15kfM4iCFnrb4THP16kehs/2p1NXL5
lRfsnz4p5mOh2IJb+moOX3cUuPwKu+qJanrg+hnETgb7A8Dntw7BqbD8ZgtvXmb2tPgRWiFoNJIz
oV5U4Ui005vAuphkRTKKC1xHsnaVhiuSQBKa056Dyk3c7kFbnDhpuF3zkQ+azbg3yqVv19RAKC0g
jvXqCf6PuJybfWmJXvbbwXJwxxiuKfNruo/kF/j99v5qnILPDcBU/vmz6mKbOXa21a6oEUv5Mbky
Ev1JX4sOUw2gcOzdB5Cm1JdZvsUUBYo0k8SIUvY5ZGSSLZWhEUsX0nAe5+r0nVV7r/DpCjk3ltQU
yd7MVOat2sCsyKBOqkPwbMajhVn1eJBZ+Kuosk7hXPbDdwQffvbzxbk1IEWHrD/1ifq7L7RR/uy0
xnhezWRMuVKzY8tLjFFj5StHj+Aauuwm2wDJyajMnRiGKogZAyS5S0/UXH7a7fLzC9o8j+3/D/kO
pu67OkXv69q3ztXm6a3+seXwc1nTY6EfEHFunKFBS1lzF+ZL/bNA+Lw4bjh7jt+jiRf9NIWlaJeE
rX9RlWRML0swJOsiRTjWNe74IZvhiklA8zJzttvbBOUMF0U9YRD0SIXgfLGp9oHjPGD1h8LVPzPK
dS/56nNmMvVHKiHNrVzhXvxgGAWeTY+MVRMW1EC+aTv0lXw1kGkKGwOucT2DVGJq+Jge/LUvRITF
Rp2Ha2PDfpqTHHcBRHdwg7ufJSj00kMmAz3l8OlRSl/RBDYkSoIjuhmJ9Y/M7gmDclnQ2zJM23gl
X7jv0rCvfDY2+7cKuJo2HG2uGrd9qiTtpmgmeo5+hK/kKkoADo6LvSLr2gyMjf/ayzyBbWPP55vc
W074GVe0luJpYbw593BHoO6wpPa5cbgSUzRriRithd+kHn9wWPGgUs/+vd05jp378LBIURLgpfZd
LjquF96hHoXAMycfMfBecWeAdt0UVcG2yQTVfPG9l8yAxTnWv+bm48/rCby1xnZEtvCH0KdSpKoC
8T0ckRCmSxtO+xBUTVcMKq7nRPmSRBGwHdJkv1Y6xZDUzzc9s1JTWkyyP8Dcv0YhUfPzXnyERvq3
I2gGcul7FpD4K+2U8yIl/Utb3DfLdKlkSyoE/L4QOqe2IcJojRGo1yZNKslJ7cSoaPDa8Ji7wVG5
a6Edv6p+cEALHyp9LBOFlLrOPj93cfloAVCrtyfPXZHbCk6FCaBAVdFDf9QWxsraxcDzd3ycyD+k
xsXsUiEqGcH6/W4WQWmB4xgmXb7x/iEbHv0NHDttMWUhYMjRCgYNzu/+6AG94Sx/o0UN0ivZnLdj
6HYO244mZ9GouACRGDksrJvuLw1MJwuaEdw630GzuTpg/015fhG0I+tB8M+YAcvuPdqtzcirH5P8
2TPvbS6w8MglCpQLOKD908tW2Z0b/iQj9v1MsLZSObv7zWi/fnVw3Ss3/L33zTHgHup8VFWMukYO
6BY4XsMBYdLxcmBJDKkmM/wMC2YeWCJ8Tizb0sjkqas9VLmvyS4aIyHyJs9t2RnXptLzISpv9xQg
de2KN94gY+PRNrIvs8ERwotnv+MvT0yYsEB8s+MbSOj17N1r5soIWoOoztWWFkaAaLW0bSoO7RZk
ya8JufnbrKgmiVrL0vlMMtuKrvGb6gEEEzMR/ljgYTTa3F1uht6UPXZX65+1l/2L0Y4BpjcHr6cj
040eoGLvXCJkIisg3e2jYKId5MGl/Z6fT1Aj2gJg7fDEiZyXxmgB7u7p4zCLq9EihwVVzPVwTrAe
KvVZE95XjZDU7+BXjYkUpEmZXed4OK/TKiE/jpgIpUG1bF1U7XDPWjmLWN7Xab/c8JDGhD4anTEO
OUwNZuc0tPNOf9TyQ9/2D+oea68xorPDGFHmZbJ1PzM1WYbGnnIKF/NZWZoAYDE/nOZJauKaZtDw
jdcAB7/aNHesn6hJmI9Kxuj6IRCjI1q1nzDTXhdkD3uYVmqFktompq4591zPED8tlu4+BD6dVAeP
KnV9c12xz7fPDXjc3GNFy09uKFw5A33MRrbIiiaXgA1RUsjr3rmnL9mqI90FlNW3uWdakYlOMjJn
CGOAW1qOCHl97PdC+utfFLS8/Y5xPQXVcs7+9fFiP1C9vc6Ol0AKc1ZhyAA3x+jqWs6zYGjcZjMS
6Q7VAOx1hajWjSlAZ4VefvH/fczkoVTOwxvOavbbO0D6Pucf4wrdtV7mWsPjsWtPtuXCMaKP86ze
iXnYET8zux6GwSD0vTRHSrwSyyv8CUKNl1Rtf43dy0y8+Ybh346XQWQYykxoX+w8acpAJJZEKVi4
DnCY0saBkDwMHh5YQvgoydnQXledj2844niJSp+93TsDl9Z+ei8O+p0PqnNL4YoVE6ZSdNjHtyYq
chN9jm4XuuJiDHjM/4W4+hfQAMrSFTqrMXQpcpgOqg2DOZyPPdbxpYh40SojRRPalZaVV4j0FRpM
gIW5uKLdPKUtDu100crLl7BHjGdxus0YhWCStSyE8k8jcV8AwHQhhxrRoHfvjccHiKoX1g/Ofr8G
ESM64XAMGFGC7n0axDxlIyhfs0hdqcsAYKVp+LipOlxRxbyCYfeWkeFLlcbKzZ5mCsyWfyIYd+af
DFbVtYfmLCXOtxv/U4yiHb8i2r4VdDJ87cMXJ0zQzyGtmZFRBmDVzxe2tFm5+jUxUXsantacRm6D
qeBRclEZ5taQksenjDxD/sy2EfUveZhYhBZ+jYXCDwav+dxO9yPgicRm/THxB5ByyJhOysHNSDC9
zmIXs5669qqAL88J4RQB5dANZ6znWfUC/zL3EIW+1cFic3AU2NztZ1l3wz5D5j+YuhjNvGLSe31I
2SxFmco9RZeSlDejL3Ej+GOKzSTK8GkRj1Mc6sGqMFSrDjQ9TST6mc0SL7u6DHbF5wzUhJPRgyQL
8GGEEGU3PM1aJn87xN0c7vkjmNyPBDnG19ebD9kCJUuv/O3i8xoSu8i1BDk4hkC6QWMkgRH5lCR4
g+nr2YpiVLTRg2ditB8tzYsdxZKf9N1/+LKLqGM9WIIK8XtZDtVYVw0XHMIZLxg7y6Q4QHwb9dpf
nH9UDiNndbUKgd8G99+HZpbjXVM2TQBqgRQYaAC4u+P4uadA08iTjSKIf582dcoDB2D2MoY/juW4
/gJTNeWkyJSQgRm/CKMkIXyY6ka7BqYziYVoJG0dGxvPaoKPoOxwdGHaI/V2xtyMaE35p1CvOFmQ
GbJMTYz48Ylcw2wUGNd7gNJ2Su4IKvK+wQFVTLGREQYwjbY4AdjnfJFvhILkg3X7kkpaZ6RDB7NA
dEmbjD2SvMJY31NNR6mSTn0GfP6B0b1U6zqkW+t1/JP5WwcKOBwGhchs9g9zsNGyzJcAc/QRZ971
uCSGF6fzswET0w7flpBaWXqAMJ6L/wKbjfxMQ5x1BL1qQvLJ0O/gHZi2aqFXDQZwMC72YpMoq4wT
UqeS3oVlXIfUrf2/1bSD1OYSedhHQTfJPMR6E706KauDD9f98AjewVk+A65rYHAtpl4TVz87LzOX
AgU0GX8ybv5Y941VvqpgEyfebAdp/cfmvJ+0Rx3p1Dv0FSvkLe4qMP43kCNJvPxvrt+wfj2F4PzA
v/yS075RDttA0yf3NiOhSIf56wiP0Us8AmTyBl+2Iq3bAt/VtV782AljF3VHiKDTvUHTRiVf4Qlq
KCMEaDDTjcbdwSAGgCmzShq7MDChIuXZ/9jWBhxDsmV5wHifdjnA/m1qAi0VrTuVjLAlYvCN4jo6
Zn8BwyfNOOH7q1MjwE7ZtFCLBRMTz4KXjnm+90T0GQoXCr5ulW0NGIAeQO1M2wgq/EJaub0JaVum
nXBUHBNrN1JEYXdxra5mg81cXZLjOkhlZqFSrWtfVEeoaTS7LNk1KsVDR665gaG02UWR5v1TGS+2
qVVxVhtJelFOHQs0HT93zXUhyi8PH5hFEhECZdjnN75LN8nlT7yYBfc0xx6EzIXWHsfmKa4BULUM
mbAl7+Hc9uAxyqM6JriVduYvsiCyMyZZ/24gqMJMZcgje0jKtNbDo9hUxn2nv+Tnj5yAF1KkMZgP
RVMhPrHjeF/BIxlsQ0gyGd3XPGYvBUE1boc6pJNGcX3rp87XjtyUjg/JPC8SqUi5TQuiGKRpI5Hq
H6rFopIJWEPHs74HDM/sMw4yh6qoPgtwQToLWzPgqllcAxbeYpUGR2wR9dpT0/Njn8Kk1dNSSIvp
taxM2OTWYdJvR5I1Wcy/87CSvvMmvdSAUOEIgf0BzpMgdMPbEhvTijVfYTjyURN2rhRwIJ4DHqi3
jDNSZzHef4XNlf6xzf6vu+SH87cViIN6ogbEeHDV8aG2xpEG/pwQQS6s8eWTNCvZIbycMEi2DYN7
J+HDtl0j6aHRWbgM0cYqgmGuazgENLUNxAFJbHtXzKCUvuQfpcGuL1EEttEhkyct8bVN8BN11dNi
/G2lkeucUQweXEjgNkbcr94+/TJxjYdXq2/Ra68z/4ES+WDBHF7C6ogYxubwHsvELQBFva38xH9t
x1CVs5YtsGJErwtuTwEuKop9ZdRHysqb0KNn5sueJ3kt5yIPt2A/ZkIVJgp+m92A9tQCJWl24bPk
lSLkqPzuFxcqI3/MglRyZ1LklK44GcTcu8JYswEb8ogLaAn1uj+UadPLBcpJf85QaH8OuYKfwPKC
cB4gl4GkiVodqCch2HeT0LtMTwav4S6X3O/KaDc2KjDnz8Zi6lyukJ6JSQDoOXAF49+Yp+pj+L07
uc0uMIOKnwFOMdfnQQ6b0xzEOXBndF8sarwgoTsNbrViBuLZvbYDIn8n57tAFTsl1JRsc+zfgPwU
n/VBkzaHBUtkghpJbLNYGf43rGTnPXDnoUIgUHQ8MhxxFGSO82Ex6HyRCGIebCoUwBgWxrh0W61I
nBd58GnftJwNFCFweyk2xMigGGhR/DD3lzBkAo7stmt9phfJUOzVZ5/lSK0jiIQkEImr6oiK4H0k
TWb0o+3EW+n6Un/jR39JNbOaPkPOF7LiBFn9NOx1srg247i+EbsuZCEsmwNHRkBYdKa+mE0fdE6P
iV1lBufYm7F5L+MbW+liZ90S6/7kZBPtQ4bY0fIVcSFu3Ik0blftPgiTSGJRyV00gATkQftRAr81
raAxRkgDiZM1MRgTqT22lWWs7AXE83wWQofabLscTPv9KBJRZJ2Yedwqj9LWAazLHyW3TNistwen
5ArwdUTK3W6lWAReI2m0sYHtimDN2AI6Y/3XA+oCu3RjcgqRu7Rrr9H2oX/FIiW5T94Ls3qRvt0g
z5s/CmWxU5MFqFAoLPA8hP7pBbNl0GnlAVRQ+y35zw8q5pzWRbIsSuHm829QIdq1dtMuwnQszOiO
+jWjBxfCyAdnB/KtyYwPzKP76q18+yYl7wUfm563/1p9HUQqJb/veLt5lN1rM3SrdPKcyOT7r0rS
gNYij+GEfs5uyNllgYAgculmUDn22jdPTQObiwDl1m36+DGARvqFoXq6wTy5yjTWQpCApmL1C9BK
swrH7LYewMB6pNTY29pBxbwSkeQo37IjKw4toh8TpvSXfEIuZqNA4tJS1xRs2UvaVIGBhqyDzOpF
T/A7hVfiA7rjVSNROJKjiOBzsMJjGXlHqa6QnH9YfzsVgwJU6TflKM6EwVFwdj8lDZN+ms5USwO1
y4nsc9+TRdMfQIgqmLdKdaewYpjoyYm0dfmvK98q+LYQAWASHBIEt9sktTrgEA6F0KUHLEvzirxY
cKR5/YLkkRvfsvzy1nVlIECkONPt/HNRO4pTD5/Qq32pybv1n7MbJbXn2PL2NBItvp1CF8uX1UL7
ZRwQPpvawfhhYUXhvcAo7WWNz7FiNDzTsJ6D5Sqr/d5DpINJh4h7OAi1EskvU3dpLgJepd8Vjnv3
/woidRriz9ZED0bYhjGFQhZBxCu9JDVTpndrsIDcLa9I24O+NVkZvpn/IPitbfAzu3KlBWW4w2R6
lmIciLqClC0R1s9Vcerhq3lC3WyZxkwWAv27tXwM2LQwoQzAP1G2lbNADbFEdHjyAEOh9J6lJQNi
AmbLSixNSpdFLvqKJhOZ2Wir14/lcbYItclwXqVqhG/s6bzxMpsiioh2kfCcnNAiXsMqG8nbnVq9
MoX9nTY/sK9wJQ8L6kxATHlljFhrO5bneTDwXECoLnNPuZWl2ZcKSCdgHc6GOh8M6znvbVbYTXCV
l9tJNmNelDWU28K+WLuJgvXhgdSqk20nZoXeDPsXFk4YvDu6uOizvZLl3JQ3igPwuSL0msdlfIKC
T1K5JXJMzSDb9aTKVC34UiG5fY6a5bmuesZMX1CUVdZwHWYCcg/DjM7OeR1j10QF2hWbC7n90CVo
0YWILfMVOD7LaUlE0KMx3jfi5SYRuOCwZlCILiivQLUlb5i12y40z2In4WWJIj8lUIvmYE8MLPxf
LCpS42TnTx9Js3bkySH4/tNBsP43AMzGKzOiDWwbRXkJGLpZ7OX0tdUlr+PNoH9qsUoikoJMU2zO
chfi9P1Fqdfv7MlAx/2FCshvFt06ymCs0vhmLSPCbRB9bVnD3LHgjgQUpXRN9s6eIC+VaXjpuNgZ
kqUGnoRMHuJeKoEGq3XivVs4JJAL6grsOMfeZ7jPpfSPISGO6Gg8bUPm5Ac9wg/PrXbi8shSXfs+
bcUbQfj9unkmvQFqW2CgD14bJi2+sWkMlHr8Rndv8GphaDCuGPUi/vsmXYDloe0KOtDOLOABCB26
tIq29BQ56pp8WdITMGzgof6M22xuh4mSOs50ctyQWjgYSGZbBbWizyTQRpsewdqb/YzwNTXBFADR
6EPeqsgcG45S0g0Mgr0Ulm8+cgJRJECSvffhmFDkOqtNz+zhCcSlshQJE0eQKBi3tMMmSBVgcWFx
ivvbDnDkGAdNDzLHY6XSDBnkUncRU/sMEwRSDaXteaFol9t1puRHFN0gbd7sjjfRf0J+dRWxFPum
KNOCg4xnSIAALTR62fZNwTPQlv5mRhHvEeSOG8TXrGgBjcdyMDOKlMEwVZORSxbkP6gHSNxpnSmA
USlc9lFPOp9TU64TYV3r2xaswdZyXWGfDa39m2wt5pF/7qczp2p3FStYhnjQRSE8Wvg/2u9RCbai
+LUpkoNNUyLVF6a2ery4iU2Xq2ocrVGI89jS59Rku/4MRtrT+7Ej8Hh4+nl5wvr8R37PknPsB5/R
gycNz3/Q/fIFJJnRTAcSb+JhapKbvClMKlKxhU9dN1x35cac/fxHYt1u+RItg6oBfNjVexlDQh0v
RMDumY4qnsv0pqLSLWHkliLYan8NNLm2qJ0VixPoKkwc2880foupsPyIBF6rhFD1uLnL3ex0xegN
8x7Jz+whZWoq4wm61D0PbTVIeoktr3nh36TINHaP4UcpOY5n8NNK63oBr3FBcQH492MswCZrvlkF
gQDFmn4G9ZKLiXyYHuJY1GmLiv7GRszFKHJS05OAGNNYwLKLUyHB3zx76twmxmlKlrVFLt98gWnK
MNjcY4LXuLPLWMAex3eLCxZqYONT+8zJ/luEPx+jVOMcqsE3O3/db0DDJ4pjStDuWUCwP+RPgd+V
YJOWLFSVGBVdPgMHM2bDdLTgNb/A7tcjTA5uh+2bPNq//+aR3ucjjQNvZplNvmza4kUwIZPrku/U
TdCgme+PCmUsVG+0H5lXpZS7ZFnK/FWHCkMoBQiX3vmgmtqsXcMLwOeA6NeE2udricERh4FBlpJQ
I+gM4DlbHBAGUqaS9kbzuvP1Qg5dwf+cjnrrhJGB2wBGIaTNKLEyg8qxprqcQlVM60Uh7lpkZkTa
MPvUbK8k8AWeuPqE1r+f1qTPju4Cfwp8q2MNS0D/YLQRf7wY0Grj5oNYSxuKH60NjmFOua45M+OD
B9aSGYSgP/LLIMW8s6CftQydOnY3YSYUzsfCRktM0KN8fCIR9Q7R5bt/YSruQra2Gd6Kk7+oKc90
NlSxBrc+VS+93w6HIUqV0U6GMwE8pn7Jt/6dNxRWSDGkoV0qaDb18CrSC6pyTIYMb3b2JIwmfnqG
vAkgzDC4NwT4CRNl8iCnbNAbzNM8AHb/gv8WfeixAIGRQJcGIU3q8p3wrhoQcWTmGRNTXnM+0ELB
QkqL/5k/1+ykYN30SRLBEuD8kdxwz9OF1jKJ/cF7BgMpu3QjVZ4tt3zg4FRh3N8x/EheMWQbcOA0
yjjuaezINSouGbX5ZB3hEDPy/cheKoAwuig/J3C7kilf1MxLmWVOUIPLRhJFQgfDcXZZ2S7KEpZD
tv31M4NOXJa/0IWkKvMgnHfmS6HCXX1ETA4HhuIAEBBcfimN2V4//SYqtAzwL2p/A6rBbb+hEGnF
5d5sahA2wtL0UHRJCpg3KQ2oxZU9Kn4UprFo84eaYO2eBvfOv3v+k1gmSvsfk15IVTWlSW64A/8S
g7z26YFA43RzcQAEBrWZIMZRuUtHP07cHyAV1bT3q6bFxMoRYcTXxCgxcPRIicp3vSHjmYogGXR5
I6n6a7z5ZxIbNXalsq7KcYhkEWL2EDZUeuieLTIRAG93AElzbGlipG67OGFA9CMwsXmirWhNvK/R
1wCpW0n4tfK92mNQ59CLOewIglIXycIlirJfzy0ngR7XRD4b00JVvgmqmtvSwkmhmweufz6CZYDy
EShvK+BpI4wvKSDMK/7FSOs2gZsv1PQF5xBXc/UeRKyndyikafzRo8LlLC4V0TRc4w8LNAPRyYdi
Jq9x0KBdqixZLe573Y6XY7CAlr5pPCtdr2WqkuGWh+Wzj/j0ovIYfPM2R39b8j+F2ZtzTITwaqjr
/HiYm6d/7EQKa619GWsxECakP+v07g4YJhFKMfysIm02bJucFVa+KhlFTS1Fk2Z4MB7cm/nlzoUQ
agbrkSjMCfhiCyJU1Ex2CL554vjduFjS1KOE8B9SozsTYnPGjslwTZ5P4vz+sGN3855ZE1WBmUWj
pTY/kUSmeQh6KYWbCzz56O/VETBRpj+CCeTqu5cYfAeXNW4GDa8LwbdL/8VEfEqwVlZTiLH1Jwg7
v4IfIrmurhYi642f5egAaisMMuLQl2qxO5j6f4aFUaslvRwaMZ9UPRVBrKIOQNPu/4YjbfSw6ha9
kMODqoxMWtQv3UG7EcjpZVVHR4+Q969X4IRjZrvSpesJSDFZcOb+N9FjfrSsmZtlByWu+a0YekQf
1inumwYtRdrQ3zh6yZHq76MJjargmgvNO4ctQPjKOA5n6+FRYKbr4pUEffut3qTnQYImrFRhBguo
eJlesZeQp/SBN/fCdGcMyPbR3CHyqgiOeBCvskVw2ryK3hpULUcY5rT6FUd0Y9LJTaDKa/fXVeqY
3uAVF3BELx10F276ZiCRdiqJ4+4QM5B2MkBSK8b/RDM/uG2Wz1SiynPw5BGPVM2NR51t+Ag7LVEM
g3PdU3F1W158/+ADeanfYGQseCQNFBT109ZoAo1mdJA6XB1Tx8aqQLBS6CALUEMC43PFXdKpD7Ah
et48d4QIwnomujs0KzUqStJ4v8HY4gG0/MfRgurMoFJCdwsELqBqlrLFlgfEd+KbgBvB6RJHzTBi
w/gHNBkQHaPBPWqDXSyND/YTHBYdkEMeuuIlxcTc0gTyBAMLShQgzp80kdvW+jgNNqrSBpOmup3K
RPYLTYRmU4nn8KvzAkWBzZtVDjBFFnXEbWZ3gZuLXoIbL8/6+Xy0PrDW/56PRFL9kG4XgCqOY4ai
44OCXS2hQluGPDTMRl8EdRhDmsQgdKXy0yKds/Kn+w0ypnA7szRb2ia/iDAv+fDxPmF5cgu2AOoI
QeZRsdPAzKPKEIslLJJCB0g7UAIhYhqcMhw2im+9q+MWzWNiaBrKA0B4OBucfZMOfEaklCs/LoV6
W8hEIfgYBHkaDgGycGbPhnLlUGxnkM5o6V+pPbIHLWKHpyuFDlNqBJ8/ZrFVVEHPtAuFUP+EcJ9g
mN7I7kqgLqHsVVd2EpB4awSsS65ieQpErJhMn7MiA9Hw0gaVSWlmdKm7eFko9BgmbIuZQWp7HbAc
byWIGXfxjdBNJjNG6royfcGahGdK5HFqnag2mDsbPXITxMduceNykyC3ZY0pbO0duLonx/jPbZyL
dBrQ1zFMMqKjE7JuUzi6s2KPrZXOP65p5jkiFSm+b3SNDEoyYVoQoC57OKYAQyddOPQBPRX66WGV
N7eKSlOBDdNcHk8OF/rMOdg1YxLaUe6wdYkMZqzs6cdtT2QjWY6+u6+OIb+U0Vb3C+H3qHRIwM/B
sBVU20wyVVIfaRGc+IOAm2uLvqWakFXw8pU0cBXmknrqHMAJ2LMsWzyPquFJ4YpBgayYFcPaUFIi
UXu9Oehk8uytN+qFEglPtuTg7owlDsASdvE5Rt+FGt489ZZVa2rRRzrEJZp5rItNL4zwNElemgxs
Jm4QgvVqRV11oZyQiZ5uhoylN6buj2Po2fljrfejKxoLV4ytr3vrW9J17lEjkcUVxXmK553+BoLh
rR39+y3xC7tPu+M6b2WCq1ncTsHO6OscfW5BN6xfX66/TpFUpcYlHJXX6BCDOHSQcnE1y8Crljsw
wTirp9vbid9gVrjylqQTZK5dDxawJ76ceK4b0L4g7seQfS732GfyGoshz06G465v1Zp6Lxt/UTwY
l2HJz7ejK5lhiBA3cWeq3s71MSaF6g8TB3poUk/HTwfX9t9+cvveTOUclo+52jLcStQm5e1kmty5
dmIXVe4TCPnWYz+wDkKFaK6nwEmbc6rhFz0rd0SmrTKocR28BEDwpKnT1TpjYmTHmHawQAgj6pIN
azmD8cDStlc6lDC/YTslZJda2HBiYZNksjtRoP+kHjKkVgNA5qFyqpddBlVuIrJY68CVfTQxZqEG
nd7x2Dw+cF3q3V5yBisT7R5r7KK8x9g1Sms5dZLtiDntVSvrA8NMu74R8LvBtTpNqAFAy6JFcnF6
XKPW04mxm7Kw17bllZEMAO/kkTBpErYnY1hca3rjNci6P0K+yvPb945FnmEkdgWYzy/Vzukvk2Rc
Yu3fatFQtTdYO6hXlnmcpSgArW3qIIOYswLDV2fevEmr2fyRw8qwLRZe/r0se4i4OMfZcd4Fey6y
Aey8JUecKEfHcVoiKFNGiLOhWwkUyauhkAn3P0ii6A5EI3xLzQLijOwrxCZai7mQieUUFwS4vNEC
TIyq8wSkVXJZa2kM94tUp8G4U8lVY/MGS+WiqD6+MMtIAuYEp8aI9oKnCNIxkj41CVejMsXXHVD1
1I23NPxr5NgEXNAKos9mcPgOMr26X3f8V70Cb0zJiHv+/BQxOKj24++ODf2kD5cUpI0KVCL5cUkD
aExtIelLikZu8MtdPXGmfgyrKk2omijsr/OwtbOuP72HMG32y6RZ9kSMo0jKQ2vwC+b/lhnCQdsi
PBUj7BB+3AoduK1Wv32MUwqg8KqdVFZweI9aqoAd3/XCymnGVL6UYL7kJ1PPdhBGOMmFKAytFNxy
RlWMRWQYU1DLhTIOzdK7AO7EGxoXlqGge7PdUkm5I4hWyM96w3x2QPpZBFLp8rEzYd8v3seEhHAX
c2M+sHMyj5n667vmCWZYw4vCzDzICfZAtYMFy7yPRexFU/bEQsN0qYRRYLKG/lO8vUyaWn8a2zAB
b1fh+L0NI5e2ClBTIjnQANnXXGhqOjtMDRnoT9PIIX9XWhniW67m18yJZY87YZml9yrQxhcsP7wk
B31cPbUUOedtCNKnqQB07XDWdaNiGRaNtJ++eb3cT0HH65NCkhxWUxNNhTiAiuMGpKRTwpsOcA+a
oMgVtW8RVlxm205FeF4qBZJD06s7aXAWdyBqvDRYahhOTCUljj2uW/j0E9pYM4dvvdxbOmuYrcOz
cKMunDqHJ4FNJZJTCwpJF1k/5T6M5eHvzj/US4EMlG/k65ntWaiHoSamEgp0MHzVhKz1QYZHaisx
di1ri2i8N+YgwP5FcuVPLcuOa64XuDNqL5gZEptOJeROhKlK8hmOtASPQTxjroHM415fJ2FZ7LYX
lokLTXtlkvKuvtgQTBku4E62XPAwuHPHUQvac4jZNuZ4VQYlWnuycOLnYeu3dcDMU3LmkBAja/HR
O/eyeO6rR8vnZ7+8Bb640FwFAX052ECif6wBF2PmXk2kWQU0K/uSCRf87VpvBXh/ub4lBwcJu9ZL
MEVrjsZHueorvecphnDz2nQCd6+r+iTdF930kInr9Vn/8MMwV7nNZVFj1aGhOO+kdab4CWMRxh4i
t3ecioj/Ts0/iT3fOJq8WfOSZEPY1kCcFFXSWFz7YLQMQQE0W6uirWlOHp4IZYKVxlAc/edYgFSZ
fPFRxUN+5kLXoN7RDe2IVtG9FtscDZcYPEeq0ne+/OWDaUY04fzN1lPXfIY4BPrIMnwA3Q8UAlGI
sKUO6v8tOvu/EVCEbQWbd1AWCfrNeiaPhY1SqCn7X7GVLKcu/SgWHrs9dZHIT8yQ8jhbOK0t7xja
dnrqfNmb4DlOqEYpik/HZ/4cP+XevQRKYgjWRBQ27LplT6iHyNJxmCP8+2frEaPvi7l10lSuPkje
AoGVQ3uvhnwoiqKU9coH9t6EEfbACxuKD1prYxp/DIM2A8PgCnfYQk4G/+4u+GEHtQE+LqAehR0Y
y0xj74DiIrxGbT3dVXpYS5U+1+V04+itueqU0A+6DZfbpCRJIi+8sYmM+Mav+ITMyCy4zSyXrM5k
XhUH/14YF1YiUbEJsqmz4OhCNNPiimMb2yh+T///1wWAsPaIVC7tumJG1VENJjPA8Fpzzsd76BNx
4r1M5yUCgfM+0CZLkb1az9WaLRiL0Z7OacTOHGc9EkT0Uh0o8LkMFL/kzeo0FKl+hrOVDnL+YDoe
bZH+XxG5KoKujOL5bkbLhZv82i/bvtdC2+w3mNmiNAHqU27KCDgQQAJmUIiyLP3WbJeBuMbpUYHZ
E1x7cQ+3610qbaTNpI2Gn4WT5ZsPmMr/7ewLuwi4Xa6Ey98N6PrGhAuX4IS0ERS14rXkej15Ydmo
0Pm9WrlKNM1Tu/tasMJwGCS7YXs/vvNB2Dw544b6uuQom8XbsoHWdwkJi7OWn7T9KuqBZ9wZqEeA
zWPObNzbrCS2HnNX9PYzJw8QFcBjr0/AC48VslURFiX8Tdk2xyij0V2L4+fON36qQc3GbPOdOw54
aIzFXK+zyiPDuFBp8NttT4Oi8P9pHAmaSVlk7Aaag1LWXjLQBg6H4g2AmX0JbNYDyYAbIvtg2pEB
r4uL/T/OhQkM1uaheuRgNY/CiVadSc96KTHpqafQ5grlugVu61U7sf7ztvSzeMY6aXuhIv06koGA
hpSyRWy1agHi8aiz/3IZ7PClSl6Pl9MWzEv7wG1YFezw7RsSwpe/LT/WzpcHNmclHKJkh6gW77YZ
LO4YHVB5jAHRmCCeH6qyT31VbDhf6MIsR+oBSp6HKQOBcaxEZ48I5oJaG7aEkDVDcpFXnF1yEnrg
jXJZtfbxY5xJaGorQ+zXLqF5C7zYzU7cyX6Zc7FbpCkIsDZBnhTFd2o0eyVGV5rgwHU1jibzrSDk
qzkyg4o7veZOQkf84cuC3O9qYV6s1cbxH/62L0bacBhCRcxE8DZRIdqjQCoew9LA4TkxKhTYpqQi
JQCFWyd3BbuAQK0dyz1vY3x+duOdiC81kggTG0L+JR/5pUayG3ghywhUKibEU0oojqedAMhZ52j7
N2xViIqiFHwQUGBSO5oOzpy7uncv5o7lngy2ReCwevWk8gyJz9XhJvIyWKaxmNQz68DpbU4kdn+Y
j3yM5P/RipCLcPA67eY9S2g8MfZfOifRZOIiW3DgF/ROBapLG0EEadrkYEDdyGydu3pcpzysrHNJ
C0GDJDJH4fjxZbgX126HnO8fOKlFiSo0fSm5QbZp67lT33kjy8O4S3wlQCcQk7rAB9otKAGrQRPp
1RpFxxYTnEeDC5NEwBwG19EvEnNdUxVmkV95fRVTNgnJggJY95R+A+hhqLeBDqc+gMyiIVf9xTbY
aO39oFezRXoR5Ag2JnEkx/iSC1bp6QmX52BNg+y0J80pd1bIHr/2fPzGZLNGQzP9Xh51onPRA+95
MHfT6EUn+YuW5dTd7RocpDMlXwFvd1b38a4pCOaeitJmPxTqfKnAf8vOxa4PFcmS1T2Fj6lLKD8G
tLx0JQoEIuSh6R9Mvjh1uUSL0qPeWfXqPXowjuUWV2yPKLg2940ItF4+EC0fK9pf13U0k1zyioyw
P7v3yB65ZIBHxWLvOweS8keZlQtvsWGjVr+BVs0WPR30dU75V3FbA/3cVMFp2atUbw7kQ2hwTmJs
qa191ymRGN1RmLlZgYPazxBPyVTcQjbpGbTs60Fmj87w0zxReUuv4GmIdp78/TBsVy2smzaUu6Pt
hRutJHmWFCOih592pTkH1LZ+saaTsmOKLzyVny/4qHobZeGtyMrxtqjmRNepFWzf/7uqx2il+Hhp
kx3VxMUwyLqwuV3ysy1Z1VtH/VwOyAFzewcA4nPPeuI/Ghi+2xJP78/rXBVG8qql9XeKrWl6pw5T
tVqMXCGdB3bb1EC7z9aTleZMdc1TxG2VyNDIomduNvtIA3f7BlZCBp7dhW87Eze/zrwj55PFPNYT
e0FNtQM++2uHaYcp1/H/4sNICfL8mFQ5yPGqCYIuxTJ9edchdknADEXgoc3oWXVdHN0G5/OSLoK7
e0fOGeSf6xs0ovqt7QcaK6qz9GrK7u2KUWrXmzbYd0bzyiUSh+qjejo+X8r9cTS7yuwp/r2aVDcm
DW3al0bzcPKkScf2S8+LH1asWgKV9GkP1uA5h6d22jc6COrYLfnVOju0t9TtdfdLP2Tvlu+mI0IH
sOu5SOu+XgAZ1UkeSRbYQWt1jL/JRJ+Y1Qgrpb042RkXjqMHYrZ+QVC1HPI7e2I/LjNW6+YzCf0c
IjM0iIvIryqzLBXUT3e2ZcT4T6aiFa+FQeWJsbd3rLlDpDT5VbD3tIoIBwHbWawA9WZbpuPZYjTD
HMhEcX8HHxIiwM336m+I3tG8nlQdcp2xgNm8kQCz2tn19WUD3IpWFazxuD2wbJMVgK5hWH8INM+s
q4iHi5hiwhu/Xs3YC1hX+6nlzXwr72kO0LqdTnMkCo9AfdUyWUlQtaOH2vangRtWbqDJHOpZB1ue
QxIUkcEW+LVWn2i/11xhrAIBOSTisf3Xbr5B5VvsSZMZX/2rSpwmK/dkoMB/1EBe4XpSZcP/1NXr
QJ/rCh9H1X+B68XIS+5JDmtwEZN2rGmDpn3ipIFvVM0MF4WGiW0OBbu56d1EIZnpDKhUFbgE/ijQ
m5akg2Zxxlr7mHk4skos1NgX9m5Ii+8tKJh84r6RP/VjyFRowkjfulg162lcaWvxZg2Xbf1lmuqv
EvQBFV/SOl9HItnGkq1OskxQA0no9R8t4egjt5O36LWBV73Wv605vi1lZkgS0f+sBzdlDvZtORCc
/QF6TwPCtvimYR8UdPoYqlzva3SjQltZThg1l66lp9BUZbs1NLu+Fhc+qpnPPWwqdjjtgDyEY38z
EzM4ZLbYhVCOj94lpqHee7knTkCRAN1dSKF+HvX8R7DstSUG3ZpgtjiDUqD77NIuIpXpxVxLyWS2
fgKnz6MryKsH0k2BveDZ0mWZYZhPIvsKdXA0Stmu8HFcTjfwcskTyc78aYlDKVVAQ+wYGmo5NP1g
n/g+WIv+UxauFf8UaCNnT1uBMZxKvjvCQSe0dG9+Xkx9Nnlo8d0WyzZxDH2dAzk4Oe9OuO6Z5g7H
sx1uW7CVnYBQVDQ+LktAI1CIckvgLzGTTldAcvdF5WGGE2chwQNTxhemDIODlRefTaPuUHzgeXe2
dHqlH6JWawDWZKGgZCkBcKUSKFY1BAjjMuOXjzaXso4XpRNJwr9v9s0PrWEZx0KdkDwQg66Jjsnt
h0DeKYgq2QoxyAapy3xkfnedVVeAQWp9cFN5wqFv4pV0fd/tbMytn+N2MTSIUqwSbWuJF2DWiJgf
U6Rvn1pDlUWJq1XVfghKSND2RyPyFhLSvtUw5A0Ef0KrrolR3kFADdBCPym65r78dXA+sTYC1Fc/
zZrIGyKmYBG/4fOwLlUVuz1mPXbp5PAmIG0FCQr1HzB6T3RKgz9to7TJpdcsm7l5Hvd/GElrWk1E
SD+tl+ZeqTKPfJfsSeIw1UNd9Lgxya3l1Td6vX8Vo4fA7aJ1rrCuswCj1kStyKuPV9HVCW3ayTP2
YtlVd+/JH3lH3Og+gMS+5caU8Ba6bZHf7XsNl6XbvE5HqTTGZAqg3SPmTjuLnfY8NwRjY6wFN1OL
/NaZryiFYgto5CRPX9ordb6ZEGHCRZCvxa4lsBNU8oZQBcD5kD5iPgDFFrOz+zMIP+i4+iEke8uR
gQQpXRSm0xze1Js7PgmruZgQQE7XP5lDHObRowXQRM0PB/eIqNTQNfnFablKWLeKSkikpKyUGWEu
EVAMYU5Mqw144ab8gkMBh5ESxHFyJtpYgPSHdYJyjVyccRa/L6xZtUNVoTrF4I2kiPUrvAXJiWgZ
1JA+NB5KzW+GqT2edxTelNLhgcx/NJz261LypZg+y0HEb2WXMfknp6iX9+4wROBKXJSO205hCnY9
WVhtqDlsgtpO4dWoC06mzusQNhjtH7f4s2kXtCLcXGLJ2FqWTiRw+k4qgNX/3qgrhh6Idzjmrlix
cxLJoSbrJL6LbU/gqQ4wwfVl7AZVTDF0BxzRl6lkZPt+SQ52bq/i6fpG/kFB8nxNMs+MdH8mkfEx
Mcf1G53Omm6WPD0lY2v2epxbME2mZ7S6njumnrM0OciA4yclqVNNl5z/yikfXFcKLdgASMJ+ULTx
jd0VKz7i6PE6U46xYtYqIL3/1qvfBQLV6tEEK0yYBX6NjW9WP8Kkx/AorekK+hoYSu3o7xWUAh/y
P7qNttqTCEwJwt4f+7RXetlRBWWKtOdGhHsLYMQE+AAMMgBLU5PQR7Nm5nuEI5cYFQHzAkUxPPl8
KUlHV9CMwhQz2TVtzzw+OYk2sE/ASWeBdPVLztEL+hK7AqbGihmwjZLTvBdC1mypJxiht5eEKSTD
axwX1Ybd/CvDwEVsb9yVWfRnkdZ2BB2xqyl6MC2dkUD+dAC0SBwJS6vVCaTJOLuc5j5K/DxVuGfG
mXYj/pUFUI4Z7SysqR9/sLkbeXiZ1IK7tRXtUsy+GWwEAdI4T1lQi+iwKrV4MRJzTocGXUhsZynV
HPZJkHul+GDcYB21GRr/EIwbxbaRXPq4EImYqnyKXFtA5imj8wsFLUpwbxY+zhhnH/unpXrQ18tP
HUlpOgEPDFWehoR/nXVkCB6gMJiYKFTITsxl0a9pYM7SFSv0/fDuoxC7YqVPY1Tyjcg2GgtBPDFO
UcmaQiToRRFKRogMX8bCpse+se2GP3bkhmTh3p1q/xB0jJLH3aMwmF3aHm47grdYzwC1CF7nvovN
fyMEgzkYLAxxKB/8/mFIjCT7pD8Tz96cxKBy4pauQvBTd7k4oFCFiZT62S/5+P4ARxM5zAouoySC
MScxO/viiFoQJgMEWCIePYNBRE4AvTUp2Jxm61ty9knt+rCGTcAFbQc0dsTW/VrmEr75KGK2ij18
uCY9aVjv9HyM+NJdbqcVlExW+LkGiKulXRPvnBZ0XQwzt7RRQ1uc2le1L/lRVSkqQQFuiqZ8YuL5
/dlec/cFuZH3J/H2POO813ibGy9IxpH2FVtRHC4VhZVeZRcEGbwi/0CV/dxm1lKpbwY+YQBOPd4L
2h6cvl1QlTgUv5SCPPpxZ4n5O+U7Fd0N9bkQgT/IIxpBrR225G25dkx2w5UDfTpQdTRPTrucAUqv
vurL+fbRsmKm21fLu2OLvbjnXI36WkPTFDCrgCXJwbBFwzcFI1Lkp/hFJPfwxEw4+3lmqT45+ZzR
oWu8tPH2awY3JYJlnza/o2FYdh/UGNKnMdKFMJyIbOZXkLYmTQDOdAINQKPP8D8/FhRGX9scqIlS
EGec5llIRkn4f+rbhZJAArEHF8LVOG5WulwRpiYYX89KjGL9UUDnGNUmggH1QAGryWB7yn4p0PMg
uRbZb800bBBsMVY+lqvaWiEM4errmwR+OxzmLIj+PU/ylbZLOvkcv+xln9by7d+uG/oKJX1g5Jt1
gKxfLyfREZJKstR7OKIlEtnggqeZtXzBkIKKixrZvFeQwFNVaYPUt96Ph8hlP45ZRs5oB64cEg95
q5XD53lWh3U+Zx32dc7q92loiMgS0NPf9USY/CavGqTmdyx6BxyEnqwiYD0KyxKFyL69xXai+OUm
ceeKBZdYyr6F1wJpcmSr1ttFOauJihrq6GwBSei2VaHr9Mxsdq96IucQ+s2AX2RTmuqOhV9iETW8
rfVFo5vt4A407GoY2kshGs5qLLtSFQGv/y/c4zDpCXoewBSBbneeJkS6BkD9+TQARGzHJMYTVnUA
xBITvEBY51kQkZ53fxzxDr3bcpcLd5wiSfgd6JfUb7dnBGZ4fh0HCBosss6x+zaTNBd6FRPUHBAi
vJWwOE2PNbxiJPUdyjnNgp/ixx7RFB/G8+gOSnaLd517ubk+hYkPPubrQrPlJqXgVQAYd4tE/5N7
7XaX6Uv8i35uRFjlXaUZfll4XWh0vDnmmvOlw7/ut5jKUNRD0RJrYRonWxDVYbgwtKFkSCEGWG7U
pxvVtzZiIQk4/XnS7rGSWJQ9cPRHKqfD8ET3jH827ASsDMk4QnGhjH2HOdrwqn+euBbYNt4YbzN1
VPpj78W0dqYyTqpkZb+Sd/RHrRFYk2eax/pwj1z74Ic+jo4YxI/ri8D/CLAd4SUppTtisFP29c9l
VozWoCClU+crsEOk+o7s8jOwcOno1YWWdlxe7+s3pFcTDhBR0G13cVNdmSq1EoHpY0HpyIdSFdzV
Nkj3BjhLJY1s4FCvNABE4ldpde+D8AohM58ShfcepUn00Mu/QDO2DxG4y4UiAlwwIr7f17DbfPae
u+cjfAnjzuq25iShZBdMMGlSb1KRfXAIkkCZdPPuonEmbGdub9cr0Oxo9I1M8yVDop2fx1IulTBJ
bmIiBuuR0eWhGpqq8xBSMeGq/JIe6J8/u5/JvrERJffXdA50xPwdfGaDjDvgY+yCtFuhE8IjHxhY
WOEKc2Sbc3zV4cTYfnrYILzuYORiZrRfoNnlkvqorOMKbL1mGJweBvxokBkYnKIaueppKbLZFSA5
/e0jrUSdxjR4AABxgSXDmox8ITqen7Y9Ux7bWQy2jHCkqHy526gim1LMgzStBdkI0K9dUUhEQt5E
Rjb036BOuVycqrfbvsQzyEHNh6PuqpOUQxeV0Ub4A7adS9vZ1R/lPWEohEvJt0b4fpm4oSpFxEAm
d2DFgsTD+z74Y6e54xNMBfB2jSQa69oRErnnbszHTBiQW5Gw34Sm3k2740TawL5GMMyfrtZn253n
0NlDrbTTWAp2LpvE6+hoErY+PQ5CQShMSBFPttpqhTRKx4hViJQKQDSIjZpC2Gs5CxW56tsA2XQ5
yKR2pf9dU2ny7sSLwxPqAyKvpnBJCqauvsD8RLibl5QfgteaUVx1zMl7+o2o9SGfSCaCRCb7Zqgq
SmS3IcP9uWLjhv8xNrBnMSGWBcztoxaUlc/I+1HpjbD5iMSN7JFlRkuHzbGhAhkAJbBW4E0Nk6je
idlmFyPlsNqtxRbFIb/kmWYLcE7bbapsGWQqu8xyfq+OOhU0qcO2DvQ4vNicrNTnrL9h2uHWMSxW
McP4gqKqp7WSzt1hSn2/WY2TUqZdKxbR4mPaJvN7+e3UybwIi3mLv4NgJMFUbFi4SnxJDS3+bCT6
2xsnyQaDwJDyzTH7qcmXDihMec1kxD4dxWNB6HVlHgw+m70HgHeSfCwuI5NLS5QJbUWEz04cawPY
CknW8xgj/dj0BaflguUzC/KL6xdI/f9epMr4zKxoCA4nSFQs9paRj+3u/+bX9kXVN90NpYniq3yS
FfZosdrd5Cs5oMumaN2ukVK1ufbAqg8OaZunlWgH/fEgTOFZdeqyfOhu8zJDcRYqW/VQqhG9VHTM
A8dl/dXmLB2Tl46kBRtTzXaY358sEUi7+wJ2UAe6eb9UGnrFxINcTX562iMwH/OzVfl5ZGkNm3Kb
nefOIbF4JzGyIBNIsL5vBf3RCBdhLKs2vLzMT5ko+fwp00qQfEix03s4Gt7uIiqg+HX2J6b8e85X
FtuFAQEjsA5pwnmsK69CGnGoZjo1Z+DGObymJFxCjHfs4IVvWcpGwar8uWEJgAyRp6D44n1VOfZ/
wr/1/dJXE4pblXY36IFCVo6nz4ZECB9qn4/D8g1CPSXttwAYfCEpRxPqELQc2SmGXC8H6OKeD2+D
vyeU5b3LMc2WNGMriO+GwEWlvNOsIV+LNQWHdqoPpl+lbT+fCsWgXR1Q+RVH/JTEmD+h8bG3WCHx
guLxJc2SjjXLcm8firWmqC12uuIIiTk91cFz9v7mWXM2dkD/7Kybh3nnQ2KGOnpzorafsQxuRAp5
kNhPlrP4ULWXuK/wXR+xa8qVLN9Vgqzx8qLd99IPf3B6nRaxCaAEtQ1BPEcTYscc4O8rYIvY9EzW
ccQooCGFaqeig9tkaMLAbbYQkLChk2gCOtHLviH5iEF8CDrlB87AKkGo74tMIY73b7IULRxOoddM
DgIKWNtFeY1ceZgtl9gfx/Gsij78D8tqGKHM62vVi9ZISMZlrE2dGIVcqMwtuoWYxQrq196ynb+y
FN0B20gG6/0+ylc44+11WpJ+6KOdV/ZJvdJEGg1OIwWfw5Xlz+bx24tJQeR8+286i0zJWsPG7+Ik
cB2+MyhrcDv6X0IH3Z4pcvnsoAp/DNR+WKWJXwBBdfi70PmupoC+J0FPpmMF9pCIEF0/a81ogFyM
kkP1bbsYNa1ivEac+hPZyPUc7a6JFQFVOfRTa6CbfaPDuEbJYLu8/w9RuJWorU+aRNDHvNtGY0Xl
K+h5uwDyGb3lkwUvnTOpa/Ek8vHzy22uiD+4cr6oSFtNtCiX3nOloLW2wvmtB8mBtJTKJ8tB5aeS
vWi2nZAS2TURf4878KfnShs3k4obgnJdNUonRgMsCM8H6YPVn1/1Nu0/lfE9PTzVfzEER4wMTEwu
GhjjtWpIfSoUT44P2eASlrgDDggfQvL+4DAfEUVoPN2Hnl6ppI7+6IvRdNWbtqFryn6zvPe5XEwL
wDCvh8lEh82C1PXND+EY7BvA8iHM9tg4Vq3tmuI6XpA+CT5MJeMfQvnNmJ+vkoDkQQfeo8aS2i1u
MNDB9giIcP5n2oWbb7BKVx9MM/Rds8JDFXKq/PAqMhQ6JPpT7k/A8r38paD7sJjOY1puNcW9kzIF
fWW0W2qODIcQQcG4e6sg9v01ZHxuMxYFuS/BeLJez08a4By1suJDQqJizYPe8warREv6EUPo8lop
Dy3b54lFCCaxJte6oes1E92/qSv1KYrEiGLHISXLRhjkH9IyXHjUH5+5pU2llebn+rLjEOyYqk+B
K5y2XLLYyE8ngqFKPRhFx9fAJAUi40PEOzh6uJhDz/W/dhhivlO6ubFCGjHqxnWftQUk6+/6rrLl
fVDysS+8t23nK8T2Q7M5vbwc5YqXvvGWH3D+jRuz965cGePtQKl22Ayo3R8uYU+kuEXE4mW5CDx+
iaxhft1D9nRsdu/0+RNP+V/lXv1sdrtRIbIsOMjwG0suJoCx58ut5EGYEIBktuJ+Ayfo3Yydr15G
W8JnqUImHNsjV76E/esR7OU37Z2ABso4G5GZc9thvOyD855vBH7ejQVlmJxEVNacjHd5TvkHDAFZ
vXbHoSG39VW3VokRsWYwNI7BW0dZwilau1DCruY8OaeYve2GchojJjN/XFYsykcdVSScrrWW3k9F
C4ZoAtTc29Wf0qLJ73HXrixCkyFR3rHnApxx39QBIM3TU5t0N8DWDKrWOyZJwL6HrtP7LrWWIyyD
Iod0H/I/96+IMlDSk+41HO3D+pcB87ap3xK4P6yd/pCqnEV2fgi5/n6qcHqVUGD7BBRhRHR0bAbi
23gt0sL78AAL82cA82scb25zXnTLQ2T05rwkqjsqOse2y8EOdUC9I8jikw+RRORgJJynI47QN70y
b6vyP5t9jiXk1yxFOe+/zrxNE+pZOS3tz4mxfCzjpGx+ENd7Z0xpMavde8A1kMVccxccYqY1kWPU
rVj/LtVYj/839Sqw0YymvTjkuM318R0+N4I9CXJc/vaNchFchUw+XBMk4sXspMUhj7FYnrR8MGtI
Jm+1ZavBgaltd48v0P4iS/lFw1WSdUfQRE/A0RjaYjMvwo1XeH6OuBGp5V+lIAU/txKafulma31k
j6RgR0M1pbBfiUr1XAV/kSprvUYhvQXDbt+tya4Ko4PFIkr2zt8BB7VoZ3yF3fWswvGRAZm4rty8
eKikSPfgrG07Zy/2Dw1yuqawdfrRYz02xpa+WUESovqnmSnlIqgWQmfisUuq4vw4vwrL1An0eGD8
IFYjlE2cV4TUSpCwVMt27PRWrvhC1tfhhDDzFmArUrweOyVOs8bBrv+j1CLY9w07pfS8faea2mkn
8V/Omu5QsesXdqtDj2jd51Rz4HK0IqPsVGFO9e6JcvE26Sms2YzSMDqKdOJsHDs7c00njuMzg/YJ
rjL7fSH9HIbqCwm6IQ36zjyB13+iqGF3oaP3Jc+U1ofLukSYXydwlkQPsru9DoB0xPG4k4HI26B9
CQJb8pHmVwXCELh6VoFsvXDlnOGgzOfs9C0TlWPbNdKXMPSeB7JTwTY0jF+AALK4VLSBWnXAXV8W
oS+dKOH5FO0IpH0DjGN/bt9XzJ4HV9xIKvfLeKQqljfQ/MQhQWB4eYmdEkvTmnOWa11MtPvVpMKc
dQxZt06OK9QbbRcT5BTqi+OSKNtNAc77CwnkQs0mXdj7UZXKtrjMRnlkDaDGY9Ia7owKOnMHNDcV
vWF8V+TUXiFRVjnZIO7DV0HcjGHueJ8OKmFblpY0uZqkgXOLT4VrwEqcDEqqXFKqppxtj1gJh3ap
NF9ElbOj/MYnTTmIU3gIBjZwJAHXkZzaOXVzdZs09H+7uOxxBAgCByJMNVwK0/2qhzpw7pmP4FCZ
0k/fLLKIoJGmZ5xC6/v7A+M9ko5W2nhRoTkmQBgU75ZI+x9Qz7NdIsTeb1Pesngm2tb7FaJstIBt
IOvDoqMtsb5T4AFWusmMlRPVum4L/oxcCMNBRFrE1ULWZUJzOKBNql4i4u0sXKM6ysx33YwPxXhB
Z0mrapC7AT4fkZEBRGjeJ0uiBcbbCtqo0QS0PoYYDicG4u4AxlNB1nsmIVISjcxZAf7b08F7Ax0w
L6lqSl9RgfS5naR4fHnPficILmTx8lNvu4JvTF4gJ8kkyOF1eo7xoRcMOBx44l2VlTjC06LbqVCL
Y1jlfwciFYz0le3u4gkJgfWcmqRaMA6FndiGitzjAkPJlIfi20/TjeM5fXkBQ4LJzOUmcOnY6dso
RfqYYWx18ul+EvHicB24QGxlCgoxsaq1y11sVro/Q6y9daxSf5aKXRkOtXZRk0Y/xp8/2e4Sb2j7
wm6xXhJ6l6EotDqRz50KpnM69uFpaj8Toh62nLbmuqiqMxdhp0r25wHZg/wz3k9jX0tigjNJteEo
069/d7KxmfbwCgKTfo6Ql7Q+beUMYY6AvfW6NSUnZ1FE0qxVmyuOyJky3rW7OrNP3t68sRjzQpFV
2hsSekL6m10aUlZTQnAmhWr4PHb7+WuQHFWNxLrzLPtF5cr/t5CHrGA2v4VnKZ6tmRWCt3+ncdWA
/rP8XRD18U5798RRC6OzzGabXtCBiEzWWtTu2cFvli2mA5M5VbbtHQScWI8/7pE3TzTRUOH/vte2
8+FDifKNLDpApo8osFtVaM6Fz2SJz8xjKnNJPnrzqX8q4AWDkEHMyxsz8c1ppYn1AWXtFeLTGOV1
FNRaWvRIZ7To5AYmW2gRe8oBhLUfQcFQuNCpz6f4nmazjza8MyTN4bYtXjyhXvH7+kCqIkED8MBj
hnYFXpYm/7u1hRxHnflfByHWcYhehV38x3Puv6yDs51gzZdj4lPEq3k/S5E+L+xV5efgxyI32QD/
3zZAneLerEJY92lwTB3i5UMP4Y3SUZQ1MdlUzYK3btGMgEG5KfLUyS3B3p29kDOhvllkF3+2R5bP
IUcs3pV7i2DEHcB0KsMS/WB71OoGARRXrs9fF0CTn6758DqNcYsRN5xIt0qazYfs/ImpGPRGnGOZ
6R86TnAjwjHm9OLkqS2/7mIAsSqN4irljzAzsBETcB2J/vZf6XGDO7++DQGlD9c6kiSZ8XkjK7Bo
OB6JPKnq4O3khe3tkpP2BH1BTgYs/Um9+X46Le5lRFq9nkDJXirJZ2IwSnoTo77OQBEFC2oBIS8X
9YHUYChDjvBAOrat6ZlDV93cSyyY5nDmindaG6TRFjJnz6IabVmt31yPflOlIAr211LRz9EhZJaf
gOsxQNF3ffuvPKmCcABKoRH0r+Ta8GFXOlSi4P9Ts9hSEATNSfHCIXGZUeD9uMjId+ABGNvMIzYz
IGNU24W2lMzizTr1/u+l98/oYW8v8lOo8tzZxA9oe0JsbPn441F0bvBXgS/lln8kt5+vM75PXIp1
FVU8EE96MVNlKsuSEPB+0TUaz5NN1sLcy3/yTDMrRQlD7Qecp8m/qTAQZgGb1cLuZyTBRoeS1OSw
Y9QFpoGKnrz7UBUVn1Ph+PnpH41zA2HURJ1XwvPVWzexuNo/tYMLknXBIH4ZSt0vKx96ymY9ZZhp
SdN4TGMqcVJx3LWOSRyksgEtK/c1vXFOlCqZfPH3g2InWmPHaIuhMCfg1Hh5GLbsJN0FPHLuQRPg
5TRzqAh2gYemGt9adyzf3BoBe3a1R9ZFjBs+DQ1RMNNaFtqxY9F3KsUof/fJVtnPufNwRwOIAeeo
o79SxhuiMhtWjzTVVyaMzhCcKyKic1PhKtkeWOOcODA7nFSfwz+RManKEudti/q/a3PGIZ0qUD0q
rXP0+cweyV7TV4536+vNNqrQuBZHiCrjyr8Fvqv1Lr5gjPgO/18VDofMuK7kBNRoqnN0Kg+8w3qR
3l8XtmiNvgGnaXWxQMQb2ldeA7SqnG8lHJLOJwthOeOxSgzBQjqY1rWbG+iWtS0JhGQK7HOTUzor
dPJjuHa6qRAtrH7ulQupEmSxnEvtY7aFddKgP7CZiFdLJLnSm8m4p1JopjCt+43R3PNW1LxE+rLO
gG9DC5WRx804x5/hKkfY5gq03k99iTb+A90uyf6erTbLTh8imtPbCjWhGkZ5XXXMdt18HPHZMDCq
wkuxTjWcSvH6FcdmlLdyqURy8uRSIuUlWoQGBaJ5wVOJOvY2d6I+xbbr+NG1Sryv/CLNYjanUhhW
nT3xX0/swv4rbzpL8OHHtCZaXefrjj0OM03ApHXM2Zg4mej0MTKTHsGEIzRsbITryA8kw71dpD0X
N42/okMJcTKKYLAo27Q9+qBT4yrwHk8vfFFO1va6J+Hr2reaikPNF54rsySG4d31NG8iXc3sCuiM
wFP4UGGRH1f9XBe9I1NDidnLcWHV+F3JN3+UHr9rPRquesv7gIKNkEulEKOp/+efFWViSNbkTiB5
7f2RQlRf3mW8b19eJH2mkbSJknUrhvE8iPVzeYgJF16ZyzPP8EVJUXRK9RATDXcK1SK0HUWKcpkT
JQcP4jDuDQbe9UAIFXLOQm1PpqdF7zAR4ow9Zl5T85xis1qv2vXDuBbfPAFtQovqGS99sZqLpJ4G
jDIbcXjdb709IET3BGshP2UQFnjNf+/wdePwtVaYImqIr/14J7EggLE0dBPMXVt545jFF6SP0MiM
vBCjV50j8pY7uEEW3lZ5AzCCKOe8ps3Jdnvi9PsFz8Ck99kPV60cUD6V7Ip3+K/hVaDP/NjaMj6o
EFVX/0Btn8/cOUpNmeyVQGUe3q1Mr19oVXBzsVty7ZZEhPl7Sr/dXy0vuIq2QrJ0FvhtYG6KD9PS
+joUGq42hnfAcyYwPyiV0qeBzVwSlBX+M/XpeXdd/9RgvD3jhMkeK9ZJQEzvWy7Hk1ejJdIPqNeW
euiHHHIHfpx5kJWn7Kbqy8WGkPfB1DguWlYndGpmhMC+3f2z9qT4lU9BozkNqM/xWmHUYy39yX5S
ilhgGCjNAQSZRzkaFhY/et5DL+t9Hx/ABvWzZaHXszKQlP6rFUgCqrfKhyCsMHF0pgBZG7gOKNHT
gTmpIYyoJWvR8dLZpvlaGk8VIwoeb0BUJJF2dPj12MHO7peRCITXAT9v5I8LyU+X1wVeASWcewPx
2M/ptc1cPXEDe8GsP5r8YrKwgqQkCRkpuyev3X1W+07y9ace4aNPokDtT2IxMbDsxryJIGO02HES
533vvcf8mH54q3BIvAxsEtaME6w4V25pzvSFmO6Cfknp9lyX6s+xRADEwQLx5fZm3oOo/hJgI2Ns
A7AXGJZzpCZtcVNyJebeiyF00YUqeJIE2pt9933+BPH2vVkixvvurk0bAjRx5V47k6TjxCp2oMS8
7kaynfH1oagrpALbl9oG/co1xmnm/ff2vUUF577CxSnExw0WYZ22c8YgZT1dMs97YwT7lqabuNrG
qsvXYbKK7nKuFsZiVe7b/ii0YzMr50gxTxE7+Jg9WglA732ibjvUSzOWbe8D/GRrKwXCN70oCZQF
XFGkuCdV0kgaDL0IPRBad1Gqq1NDYF3yaG/8SSvcvGrlxTL4GHa7aL8anY24paxWGad+w3D/Am6a
IDWGP6OrJCfvTrs8qAdhhfXmi6XXZbCMcavttJ5Q9RLiZU+yEmAwEy5uKkEpVzCzXNVjUI+YFYig
Bl2SASDbMMgak+YT7QF+1OIpESI5x4R34JSDxYNvXGR4rosiePbjOc4ZWs45zlxXjl0EHVNKBqda
IMYzkr+O0we7lHzZ+C3BsYp64sU/XGR6+um417ImJZUYDszPP1ksQExl5aTqPqyc7dXzXjNoKBed
FA5nLKzHLY/ZvxOxbgZnT2ZDtbTQka0vNizyuUVGrMLNmR+zC1TYuWqbwxByuQQlrSzu27gp6lH+
dSzH05VhV7bU9zALjNpHRosdfC4YWqgso7Naax9NYp91OcNfzIWjBQxavflWpzJl6lZSGDx0OEPh
ZP87sddRB2Hp3q86rhAWSLEHLPbS7WeMPdmGhpWL9Jakm3FUwOtWzu1FWQN74bfPDwawnnyg5CwA
JlDNecEqYzvmaWnl3zt088RYB5MZQYq8zIkOPYAyAiKhKU/L1puNLYOHFzFVkczcnq0m7u6z7uuc
WWqIgdQFryKLAwi9dli5cNM1I3FoeHZRKUzAQlOtpy0Ocr8LlA050yv8lm6lkV6wRYFfmISCFHdQ
yvLy+HpIhPQ0aFTvenCVD9nFRwEAFlGfWb76Mrw6rdkKSbhHLDx5xxd8ss2V1548F8jWtdafHOp9
eDi4JC9wp8725JwxGOs8TBGHaUzTdPZczrLl1sM/9DwRtkiND1wFUuOwtFbNV2a8mK3hNIbXCceQ
02bkLZUHr2801OcpC6fCF5c4S2ESKpM5W3/ZHRmIRSXl8f87nqw1yTPNEveVfsKkWTHnNVN1CgQY
i+NfInUf8MWgL5he0mQ81rx6zrfs0dfaA4hv2zfATrBdPm8UNrteyy5/hEgYrPLYMgyEhYSvRvms
uHscsL2gBaYCh6p7KwEpYby9yNgW/CzYe4jrZgyYFAeXc/qOKGn5ppq50de9BTVsd8Gl3htnt/k4
LbzBDj0iuKZ542lDJE6SDBEOj5plrrstsDxmw6xFaKxOMDKp+DCTmv+d1inNo0dQY8pW3EQDJN72
jfjcz+odc/b3/JAgdKgn5rgyS/tvf4pAaFYOlP77mkBWl//rTt5KDxkDLalAQyxXQtIELYdrmYfn
lsm38echNVRAVsChgqJy1HSnk5GQETm4gw5e6UTtB/ET0fZrxVRf8vfORRpbApIM26DzLvQQnM4F
uq6lMPmH8n+Tts8NE4y/lenyo5Gmp/oYZN5eR85BdrVLqczKBJpDwNuojt/XAUztIDq5n7p9ucLu
4s5NvZDOkmwAIc8znesJvd6gzES/304tSLcpxSpzG3KceolwE8fpspRdcXVRc0YkbzFdVKTtsX+G
Jvo3BQjZ9/h/y0jA2VfsfPRTfE37rKmVJmt8hrsZLFeeFMUMFzLlA3BFjTGiQcBkdWyvGJV/DeYb
M2h87uJH3yzGIFd2PntqULi61pyCARzr2SRFl6na6+vb4hxEWG7QVpttZoJs3z8Nk8ZkWjPCB0hd
Ba95kqP2OVMFuQOxlhnb8T2r5dv9SoDmNZ8nuizbOnoqQcjbQsKoGvYyEgyAj3SxBU6j68YFVmhJ
YCrnyjPQBF8H5IBkl5weBCA7hHnQgd6uQ4JdH3TUQwJeBicsuoL572rLy95S0YqxMJ5vOvy/Wv40
wSPF3RM0kb6E76YYUwVgFo3872L3TMuuOq8PAlq5VtEyjGB93PPtGy8nh54wLlIBmOaF1fBxhC7+
xpHGhqEjMcM/NXnN9Nozxw6nyIDLSGnHdYzNekbypkXYZb6dTHI7lpuaoCFbi3+Y1LLyQA4ubOXk
ZjBZLVnzCvSh5WqNFOckb354CPwhfgLme0FG7Cv70qaMg4/k8sZzbki8WxLxsI8uJYwCmQc6/yQa
70VYRUd1lN5bcugFQEnkLjBAwrsEv5M762ki4clZADI0S8K3fIdfGqWGuPempiy4+ca6n1AB9ZLZ
KH78BwUJambIl3BtD3G1Lqc4E4qUAX0+CovILTEdT7L4ulauxVEXw3HjoT6NC3RnLSdW3rVfliez
oJm6DcXEH3qFAJycfcolKd5G4wY9Y/niacV+jE1C3LcbLRKo9fD2TTVoBmLz6zxd3+HZpvk0xQSx
YQrmpQoRD0ijTLExBhKBVYy1C12bdzplOL+cCQkMA8waQZwGBG3SVic8ZoyoMbSyruOdLepw2HKW
NgxopGQuWhzc6PZw+UG0XOIHFYfCr07IaoJhySCr5BcyP2heePIIYj1dDBktQnSrpya/+j2RWG8/
i3t/KlmfjOLSzFgl3nA+q1dCF4VHpNQ270v5UAfS8MCv18KOMvcAzNn/xBjDhZxu3RQHuFiExTWX
17yvgx2wgbqPqdyGk2xop+G27TtKjcG8UnxvltTJ6It/qYpdWAjLETzbjoXNL+4xTT0G50HRqbIE
HxA2Mza/VuuQozMkxNU+OdyhJ/+2OhBaK9zZfOKD1qq9L3Wo9bSRw6FOt6l+m92SGhvny+a/ipES
tDcPiE3kwxUqlp1WbLxP8iZOocY1e9//I381BUir20CPD+/cBBIozEAwYZVh/e+OA8s+N7ViV36k
BB9qhis5nacElWmnv0O1SXQiLK+miTdmHqse0hKwqheUPxRs2hqZeeG1IL6wbgEcYi33I8ARJJ31
7doilIf8ym2I9+U3OzwnCQWpCNRkG83C+CR/WKUl8lb+rxR42HPcyM67nInlfWsQq3BhlkhYVKax
G54GvPZdaYMDAIMjemJ+P3fn++Swts+QC5v7idT8p5w6ZaelJw4dKXcU+Qjx4QJGeQ2sxwgxxWwd
sYQ8Sv7KXiY6IOHNmmMl9jsJWXCa19rGF64XoivGDnAW1wa1mYKLUrd7kdIyGJBzLPwc6Jmn8w2D
PGXORkuuXUp2CKl3RjiibGFChyK8MeG2ph761eO1Y9oQ015zs/VB6HKJhmwsjLjKiHHCoHdDVI0e
iYKlVXI9FuKLIs6XoMMiFcy0a+kM4G17Bwmjx3ReT16ZazmeWbohDQtVhYu+izfioCy+l02lvCND
rF1HqVgSJo4JYI6Pfw/nixIHeE5TzwK9xxV3fzV/Pu3H9IkzgsAqzltDj2ykJvcHEyfa+JGgoMmg
73xge/jCAvI1utqeVELCeSBpRWzQLCKHuo3yZtY5hMylbT22gMY1/4WTHrY4SlNG3B0vYYl9cGbQ
ftoNWWwz/HcCUn/YFf4nM5cQFqHioZOZrLStui3t6NbBVcX8R2hMfI5B8Zfvh7Xt0P+jTAHPFOAo
HOkp8NSxfzf/CAgsJP/Rkrv5OvVdrnYIzI0bXjM6N2ClZOsaKb2MqCXbJjthb2k58JByIUqvUKjj
ksjVGVV4dXZJdpxFBXf5gcBEdKmAh/DvNY8zmY4/vFf+1Pk2XXa2xdBDUCRaZ+YkVQjLRJVU80oC
gPO9YcOK9n/dqG/8294lVKiihvQVGdrfMopKqiW8gOL6Av/ulDS31IQtVTHr9j5iiK4f6v3jDWPO
2+PoavIyXivbqJPbOsuVwdjp6lP9L+m5ivOn9CJDPs+QyPD4HlE65kD+yKRJ2y0HvPmVZQsBGjaa
3hzhsOhOj96DKY72wkjp6+9VbsjbCgbDzCzVuwyf1OQCG9UF0IDFth0ydq6RUgoCborq9bUubCN1
vTaT6/20cBYPHPGETLISLteEM+cMUNH3fpnSlNbygcHi3X2+4KBr2OUMDjSCbg2LL8WWXqcaXAJT
oIstH6zXx569Y9uKk4iBtRU5MPVYdd03MFlmU4rPyRfnDVoJCod+thWaoXsUyNBFhKq5UWOcgygz
y0wPsuFOIqzFKndQNX2n3CftXtO3oV+/DZVLs0nyL7FqQBvfiX2L0dCSCSd/+l8TT5fv0D2wH3XD
ldO2Dj4V3oxwvmXOv4psDskt4qUqK409ap0w1+g3r+KE+Cu7JEInTzA/H+49cX+yf4Dp16OdwGra
CIICGxq3Uv5oZAoJixWRjGxMQnDsd6hVYFB13kdVj/0wCMMD44JVUVcH7sWpm2You1kyhvYtbRyu
ih8o9ftTCgPkYJrO9J1Lc/znMVLCYGpac95jBCggJ74eOtQntxXtUaep9rWdF/liyrOB4aXx0d6L
jIrhD/i8V5wK/G3sR2Az3XgBxgXCmbxOxQnwBuxIySkHJo2KFfdMyWEhlgh47WLrHcPHwM3g3ymn
HZA4f64GqtxB84exMG2Lj0GgLeVDMDYxXioNrnEo1KK77a6UU+1ZP28ewoxd35KiC3SgHjJ9+GIy
WUWQFC1kTvDKYmn3N+K1WxZ6XyTuESZRDJ2HFm8XCrl0fQjrqst6HMWKBTdoDjrjYCkUXfj5tyxe
XpRCQCjblTuB39WwBZFH/MwekAWpANobQX77BHQ6VPIY2Du4XJEjs4FKkJazTee9rH1xMBFzMdLn
T+WqIGxO2qJaLGBcKu6e14TlDkKt7LDKNgMnox//LE99gCNNObdo/pDJLy6rXVtvUPWt9n+apzb1
KTUkTeFFuk9PiCcXsTRHs2/oS9Z/IfSZpm1sJ47aOpWoV1A1o5M0g4gABaVm0KjNF8qyVBacJl5k
aKYreLkEcZTUgm0RRfxU45fdcnpfVjByIWJrvGNij9oQpCG5ezXd/1/Rl0GQZnnu7jy+g7m+i0KC
HVWBRnOjPz6ux3QiPJJvw9Kkby5FVfzmYD0AiVNSV0J8SiUE3gG4glHrbYyficKCEbioGyZG66aF
VL5imTxX+jvJxIZeWt20/318BfYwN4jsLim0p7oQrSfQqCU7KMUbjMSO0b07c4YYWYYVKd6SXEpR
31uXgRgisfIYx7lSY9UCnAomVi0z84tMD5yki42miB6Fp4hlySKkI2nrsnCrOSliiIr+6kx6boll
qa+NEMfof8G4nzJ4vDzpC5qjEJEiZTBYdvZNyKPSz7jKEe7bHuZAVrdh241w449gAcCm2l9UBVwD
ole5pF3qvihiQAGUArIeICsKmgKdPhIDIysIa0Bg1D6Iv0MuPHKeuC/nMfjTIGJj2XUNce3ZFSgB
cmSvQIBA2tzElTwv2Ex9l+rGWDxFyA8kGjBZudxw266MmCriYY9Ae8bZOgYtI10LGmWRmoAW6SfW
bYDapA2zdI5AXxMfudk0JKElSVzciXcRa1WP/+xdz4bAzMG1Lah/jHxdp2wCqckHa/G1M+VvFGWK
zL9RuYEikblN6pHcmXpoTNcQcGD5bZ7oyYtMA9jqxrDAvhrXrh6N0fPmGD/8nLMLHFsV4qcEqKDA
IXPK58oY+GQ5tCVbzcjXMLOfBAdjnspC9M6MeqksJFmWwovj6v+F2lPvrwfrUNqjaUiZJBKI0nzl
VFlMwL+TzreroRxZO35r2MRa/HoO9C7Y8sAJ3Koi6bVJ7FoKNRncttEvAtZhZBZBAvkr5e3bw5xk
TkFQol3xR6g1j0aYRgeGRkoraje0t4uOMqQ/nIeElh94UhCVyHnBr6aKXpa48j1lUHru9rENuOZG
ROfqUN2mdW/aDRnkimxsP7bu3ONS/nVnP+wqRSPOulr4JFc5cMGAj+UcKdGsFaAIUNDg6dkJYiVY
S8jdUvkrDAJApfYjKxcQxxbTemP3UFvRpgLsspqyz7/uTCsbjlBHnhVTPS25wovWLcpOif4lgHx7
ENlALIQFzpIXXcQXjBkfQitYt1MtcFThPPlCsMNv+fiOmMhyOtfOzhmEVve/1zS+znZxYAyu3Fh8
z3UUTPcFJiTLTAJWERC/jiGzAIqkDcOH6Z5lk4m7MRkr+1/fO8uX7jnQRU6FdbHrVVy+mmJWz1cz
tiZdGbIM7ty5m0kC/ocZQLRefTnCSZzbpQmEGG40mGR1y1YehOkNmpr4ysZwSUIK0mL27tJdRPi8
i6niJfgUIDFD/4nkUqpIa83MiLahIdxUrLrokhAitv1KQZsduCa6cB3sCfTwd03wMjZyfW6rptgu
gGB/ixxDJk8XglAavauB/8l/sgYoFTD6hSSwB29Uls8GnTA8/rDL749wHmMuSa+zxwxJ8EjvxgIA
WCEqod/DVgxNsa2wWxMEy5DG9gN7dhrfiA32wlJAITelgFCSqM9nVbyA78obCNEgE4z2BnxnEJ6d
CwBmSvzbTVIV5YmScXWpOHOuZ6RRWaS1OL6aa2hLwi5jg7nyO7zKXGxFS0XKfvdh/+6h1bnQFGiI
+F3Kvd/tYuMiKEIC329NO/cWlDDzMg3TdWVibOZ1G3eOas+urXN/FdlL4Ky1xGy6d+1jATp6BCTs
aSGmbAjy6W39eFPVoW17lutrbl40O9hMy9clKMHrd5y29G8zw6dFf03/hy/lpoE8Al5q6MGtWKO+
WP2eEsFuZHw5eCz8Xc1Tku5+o00idTWxIVZtWhmA5WA1JRORUnWZIAnCpTiI2flO5isWKCqFYFW2
K1jNmYW8oz42/zagjDZxlOIqQZRdmFkxKfZfYycg4+2qXQY5KlLUTksZCUwTQ9pwcHhhSneLfviK
Uuf8zu/hyineWxecSKOcyiU3WfsX6MkamLSflmmD9sHMEpSGD1xMfDS17aaLnlx+04RsWz9NiUMj
zLxaXCVNBp6qjj+lFksTmd2PFkJzXwXbdLwLlhH6KoCyJ4UH4/dt/WZIy4CPFDR++GnaDprQAjTM
SdrYZu14KuvvUOqs1Vs8Asn7TphQoNkQNF2bqXdzs4aWODhpIfTWmkeOdZ8hDxoguOzqQm0AkdZm
nebK5hLpgWGP6pJPKWnUSUTGToBqOTXKGxObioO6LAVDe8DIp3pw+MLoIx5Gw+t6hh8i4RpeoYx3
MI9zXwnA/zbDto0+6oWh4NUQDfIXMQOyjlbpRzx4wuK6MIIBwnRLVpFNOLLQDNtX6JgVQ50SazX/
nyYFOqh+cvM+b2u6ePHeiv7iesXwYQtZ3rSveZFNrhftNWO/loh78YXt4x9nccFj8GCQxjZ/pQNk
ySdYNaNOtA0eWsNR0pi030gCgzLRSW65eZ2GMOP4GhgCWojg6EEtIfURPJR3j7bRYTbeFM36DoVS
Y9HNw+ypKW0Ho1aYy9A9ICvFq7MjV/BaHXqQw0zCUMsK+n5dR49WhrQP0x67hUwzKLD4T5Xhn9n7
9R3hYMtb4CW6r8DQw0ruEgFWu0a2SCAwGBBksdZGHYQ6o1mzRvfyiDCT+IokNjAD2lYx3cxAZQQh
cytYAA2lbMyJ7ORvmTxG2wdvrP0Hq8l02Vl0CZH/ShJT6Gk9ev2Ntey9khbFpNWHyNRA6C7itDqi
s3n4Ed9lr7DotYBhMdNGXATIYVzd59OCJNN2M8+qGfLb2zhBCMd8K70Qalfy81AwcIqNJhIZeDjr
//4dMkwbvYiHVyQD3Ef8a0j/18yLTYwNHQyx8DKuWjSm+pBv+TwiDpXa5E5IZZw9sAEeg/pS20H9
lquBAhKWL9M2RVeaCiLDR8srjpnO09sv0N307i8C3dZf39xRQ375nH89m9TCZJ9uH9gtI6At3rfL
VeVolEhqjs1SKxnASBuF1fTlWJ4/rJjQTR0oszK44zCEZjJaXY5dRULaeXBzn/sERZFgwUzFIbAv
cqu+QkbM/b0xeQu8CRizDimD7+KRGs8rUUrF9fZMDxnP7jrPrBQYBYTjPHhjvMaqyGBONoH2nQha
OoNeJ5KOEn1kOB0aKnLHuv5b3/HZw/XU1ix+ZVXdNADPpkRYu1veY4hq1jJCXmdYdlalEhAb1xbV
2OLwm9dGZ465pcVPFoNxQMpCHfCUb7KjBTyA/BNdjlDZ2rrkYKptl0wKeloXrM5n8r7TPGLH+RXD
Ek//W3qtJ+WJWaG1mbUmE8AyGYLOIIaXv+/4O3Oj2aL3DBKq3Zw99WIH+0j2069eFYXJkS4QK0JY
S+DkKcmNWmKHaCl6keSrMdEjAno5QwxWHAETEWZeMZbYI0HDy9Hfql492lsr4tNZtHlbREmRHiOG
vfNbpnphAOkfa5pkzthHEF1fTK5pCBkYGudXB0Rie237zLPsgcDowqfj5nzal6OVYnB+AMdwX/bL
MMHfUtN9yaqBKOT0FJKzSfqsGZQzyMy5hq6cgY51esxyata985DQus8vCDkTJ+GRnFWDMGaYbBqM
rLR94n4rggZGN5YW3PHuj4XK7QNnXIugBXLPYpiwtAqiIHl1sRgUEOIHzbbh3diSdKpS53//0ixp
7s8mzSTqNtcR9CLkbsCHCWa3r8q5u0VoTKUFF6alWGkY2hpplSObo3j4Xh6LAz/5KXL/oaqilXod
xz8wNnpzqC7U9c6pqBtQPxZmLFq1zlJB+EQuVaXm6t3cBen+0ZUzy+7zLEUhKoW6OtCkAI4vhPj6
yfl7PB0MsS+0/NIkLljNHAs+MWGxHvLuaDSl7h+VVj6TnFkEPYJp9ZUD7uak3lmgE4sq8UVXhw+E
TVxt2jPRl5X1OKFbR47jK9Zrd/fCcLDeMsx27bBKDEbDNtLl8e84x/kYBOdsREuzh8mNI1WVNS7X
aAubDqc5A7w4Q8bP7za3tPMbHU7hI6xzqqGex4ikKMVG0tmAGXkoHwlPlndb93MQUjfjXJV3U2JS
Mnrjy3sDTpiJZ8ZbXZ7E1ImqaVKQkdHJLb8YoAu5XeBOfHm16VvLZ9P0TN5Ui3UQnSy6WWrFFzQ0
+UvgMh9QIrDKw15Po+R+itLhTtuxXW4JClK3k1HTbReaG4IZS1m9oNGJOGHahQsWIIurCXuhYaCU
6Iah61ouAK9qUSF1PmZmYz6d3EfO+0BQG6klTrQNaHPjHwnvQawoeeUmqa0yw1rD9b+UOS3z07lg
tSWJCvok+4/k9FW2FoYj2m1nyCqI9jnqHP7bbWU3IC0+LFNsTEe1XaxlZ4Sf2i+L0MIcpdxEEXBq
6EfT+NCIFy7eFUhLp5ggD5WK0qU0m4oHYVDKQo49UJdZTRIhzI3jus8rlb+jAR2Z1StjrCGdB9uG
pe4HJ+GWl1+K8cAy7nLkPhsbZW7SQJAWSBh9hOHBuDI55nK7fkN6KVtGcIIQrzwE6fCc0ehWZgIE
7i2FUrGrjxgE8FJcWKZtshuPqpJeTCDVAVQo7y94mN2nJWifcxJhS54yMux63dK3pXtjwAV8NXjD
cDchRNqRkR3rzAP/ErfClfYYL869Gut1ax6GraHnnQIrtn0VonFq++o+5zdu8Sq+IizvivUFDWFB
386lKO+x5OhMZN6SxxUoBFD38BnUHdfzGpB3tHCCbR5y7t+D78XXXEmmnxGZyFK2NBaUCIBBw6WF
HMXbzcjnesLR5jRRh7jNnOAwKr/4n6EdYwop1/Ltro9dUbSzi1Da6jsQpshFwbiDl4qMaivhy3NC
4GZbePlee4Lk/Ayo+DVnWaU4BNjKY8Th5SnpKUbkoUj0iZq3skaaJJqxPwPUHW3chxa2TYi13gAm
ruIg8RY0LIQ45yf1xwMKGLuaRJglk1LHwmQRPqMcxAPpHqytTLzolO5sWshdn3EixuxIdhuKhryr
ef0rJa23l5pg96vGmQbUkrmwbB/3UCmwRR5UFSt6BJ6DUOD52OYpIF8rdEN+4nzksbiKQNDTlQ5n
LmrdjfspMnz8B/9jvTgynf2uggldiht6N0QgQBcgBqPlO3W7huJ2pCymQOOK2LJPSq7nXH0cFWaI
wG25iBHDJ813ADv0Aa1VQ2+HRXKMc5kezeD1JHpiXRKahTE65jlI/hc8OrqcrL9tqhWcieUsY0WH
9L1GEtkqedEFPRmBoS7BvdKCpHWbPaWNGdFHS4DuEXMD5ZDbXJVxa2o+IEc2uZVDtPDnen3EWxKz
EAUjAvf5FxZ/Y8ic7rEhgUJ8V6ztxzivo0Isie0GscpWo8R5NP4v5xbAZQTsiSn+5/aZx1KE+uEs
2h8YQC/bnqpAADZABrTcn4rhPaMuWBE9r61WeJHSXdMAA6NXEKwwPN/1rbH9qwcefK/6+0U/cCLh
9T8SkZtZNR/QlsfwgSvQF6+SoUfru5/41WFh/U21hPmZMVdM73KrhRwUQKiTrwM4n1Z1f9wQpnFS
GQHHhJr104YylWm1IIMJD9UhQYJk2NRYT1QqIVc3QkGUiXUGTKV+nOrJlhXt2vfiBoYKOs5Ogqcz
IZwYbmlGxdWj7s+UDwW+UURYd4BCleNaGQz5w8MvOalvuZiBmq1TB72Q6LWzMuj88riVJu2pBZhE
LB4pH2TtagwMNp8Fz5mmckW3slaF6NjxIKMTeyffbawoqhrhQM8P+9PgSAYWMK07Yp3DtKiEgnpR
DmfiGVqxPaawHCkHiiS5cP8ow8871vwQh9E9HoIXTNr7qmbdz/l7muLLjJdDO38cvPOE54whRw1Q
PPDAykmQOZ74Uj/p13NWgntP/loHac1dACm8IU0Iinopj5GCkKjtdXWtniiCEjrekavu9HLVfm4k
xQg6wCfGtu6YCJSrkz8mJzLbfRdEMw8hpzvwH79/AeQSQExU3a/+tVeN2NLnfJzwaAJKjoEKrudo
T/APxv9hP3EP4vTi+gSdOXZ13hgzAujGPvUWH2JhBhOaKLAPaJ1ZbUT8BAZOy4BT34z1u74Jgpqn
laUyc2ropQweKPm7dhxsLllgBV7d35uAHineKDozRhBaqoAnwFK/2/HIlqKRGrRcq2pqu+KaD2TE
1x4gTqZT+74JQvKPi20cD4HHl7vmxy8MOgy2nLcDmma7XJWF7jxbsWBxue1Xt5tMYGCIUVZmmDtc
MFRULprOMK0QBQ/SVVZXbsBoHZezP03s0tj8w3V0Jefvykuvuz1LM3DSd7W7eeeblEa9JF6DFjfW
vXd9WsPq+qX8Ppu1t/e9nrxsiO4IpKApTOlP0qkoiw5gMU1KYPFMwN2ELC8hQ+o9HVkUSquexD1q
ZAhdVABb8WSW69rMR1If3vV5Ga4ZlvpGmyxe++/q8teggkJbIp6h7y3flgDatvCwwvLdl04fGAUl
wYyXo/t2/QrqFlUYY9oNpBk+mj1vLNQ9m+VEbGe9V76pLyqcih5RbAxKiZjXhQ2F/D+T+cKe+8iX
CeMKLi/slWjeAHQzwqwon4Zhdkz8cS6DLmihQWq0W6CMRatnxuZaEniCsLglMPPhiVNvSFmJipZS
Fpc7kfgb8dCiWFzn7E+XGE5w7GLitS3J3gCZRh7IzT3zfQpYcKQ5+vYMyIG8koCr1bUNzQhNP0oC
tj6pVZrFoYC055kewkn4lZaKBvPtwi7hzpCLWFv4lfNnxvjXUMgkq/28p6tKGxxoQJYB+lMKtu3k
xVKlvQvUA6CE8+8/k/fPFq1amH5BQX0QEIzkaQ2wJmmKKMxKMOvgUB/nrjhjW4gxQhUy9Hwu2U5D
YSQmI9avX8L9ZdLC9/b9LuaUoejbfvUaFFXw28mXB3iEAhvOkl5Vtia9ZY6g15UwZa2cKO0vZHtL
TKTvqbO1KMymLxUHak13FYnTePNIUp7WD+SVxXsS4q1B1RRH6lFcSN3MCic2hM/auizfU/UAOaK/
C95ZR7085FJdwNhESHw3umIhp33Rj5558fJQGPTypudGM5AuVE4efEnjQ4zGhCxuPIDr3GSYEXga
yH8nIvcA/qRYt6BVIyk4LzUupL0riGIAuBkwKluY/5lmaUqU7NqPAgOzanbkNApHIjUI3fAAXyML
t4pITHoKJXhb49TnqSDBrWrUZ9qzj40+gunOZ8nUaphP06l2i0A8AbVRLHF0q90cxoG3Wl6sYp61
KwRJVot37I9MxLQvmb53FxnItCaQkTIXxTSzV14yaUSlIXYyRh31cTh5MqNSy7ztmcNHBEX+9Bow
bP9r+pwX+av8G5HZNJ1uYK7u3F5j3bBk3ATkceOBRCneuFEhCRc+7g5ShC6UGJcaTNHp2OE5w3cA
1UT2LjxI6zo95Koe8uYPOyI3fg4y5eGbY47PMXaImfmRUA0r6SFRJ8p9O7kyuDPRiWEnQj7pjk88
vnNYaQM9z7BzM0kXFQrkzDP+HtXWFsmqs3gJNIRmWA+vRccdjnP0hQEcauUJ9GGivY4It2fMCHwF
0hqrzievaboa41FBD/PvLok2ZMNqr54y1iev9TsPqywCGqyQj4QkfcEXghf6cnbYVeFZpLWXirxt
/X9btF7qeatBEcA66L70OZ160PGmQ0gGqwZGptlk50pdjeUKTeCKlgaIJuxNUDx6XSPMi+RZWg31
ncu4UHm+57tp1WlbOpNJiXSxib6ZhRI0hWdZMVEhw/EUqyNwpt+kql+6aOFOz0Ktz03Uhbcfvvn3
SFD5kLXoWKEzXpZnelLQuwJvS8euz/xjEMk+EwSwcESvh/RiEbQ9nzG4+jXv4iRDPZG5y2shF73v
GrSfIR1t4KC4N4MVYUoPaEW8OzhkM+9r9wSSueHTVJfRQivCSH/qCzKKmWI72qha1uDagEXZH8yN
5zDMlfVRx8iruhnvlkgY5bmotSWEgd3hcKXMi48e+ruIJw7Z8UcwmOgFRYI9zgeozJrak2ONLp30
2ifyi9ivWu6Hru9UI4ccl7qbzwPWPiq25S7HazmrcPWA+KwVdY+xFmOlvX5gi9+1nS+cPMoAYgho
sKp0PqKVGIh2vXZI5OMnPt0XOncC6b9K6GylV3qm+qXLzXVtHi0xU3YImJglfApH8ilSA+P8jxNv
0T2XXCsLRhT7TpEtVI5OKqiw8VD1+BxFTNM30tGj5nCjkVtZoFx4fmEY2FvSFfj3wAwfSW4sEWTX
BD1sXpmve3NEnuNBiwR/+RX+2S/4tE2zr2H87f84gX1TsaRTxop14cO+X+SFpXE+USkX7roXf8As
tTasvIRmqUKVhCVuzEB71qntHytVb2shgW8B37v3KWTEV3XtfONoX8nPyRGX9lB7CqY/w1ERMF0V
ZqlDRv6Antn6kbY7PS37e0sNdVxdYo3j4t4+O+X1Gx8gp+x98W4b5Iw5G7C/TREflkiyxFci4Xqo
+MT+DwqZ4wbBI9LsZvbEMX+16wd8mnnpTWf2YktVTPwV6Ip3NhSee3Hx4jsf0me221dYUNN5EhA/
n4Zi4T033kaDuotX0zA08Dv67CdxzBrdt3gOxDyJKaI5a/FT2/g8nO+Vm90nkOEEWskSKBXkYr1E
jHZ0DV1F9sidr4JjV/7EqZ0X8RtXp/tyCNVrg1oe2Zjbe1RQNK5hpJt/ICQLFOCFYEW5VTA2+sme
gATvVP+t6BimMz2BpmHBhSDHvE0fNefqdftudErmjL5JadenbJ/JOstz9RpzFhHf+rlkdY1O/lAH
hANNM8HytLvDHy+wB+blS4k9inqFBvgZExSjIiPa+CiiJdYxsGVm9IujaJ19YB5qblvIP57X/4zX
mV+wc3/cVKhPutcFYb3m6rhEAKV7OxmaTYCzeua4ifCpG6pd+6xOEXBSURP8kYfZ7YhwG0mx82TM
RNZU+sUPu1Yr+1cjqPmMbNDE4ZUtz+1TSaRf95Z620lN6aK3OCZoIhA3kOKNp2EerIhbih7mnGJV
znrGzR0uO7EGt2cW7pwDGRJwUT9qUvAvQHCiiuT+ftMoAnHCPZYwXBeartdKTNHyz7ZelQmzm3bq
XVvjyw9LJZ9xqVohcfhCX6RKP0jW3CvX0UGxWTz2UYTAtxY56svSbTZxiEua48oYY4LGaDDEr963
qkmLLiwtLZeWxmRWWIbUle74SLQhSNgC9fLEAEr3bTBZYcd9XlVJ6Cznj90nvq0zdbmhEKZEPjno
75eBXratxcn+H1LTnNbDvDEEZ880Q0Ey8uG/PFuVNgiviOn8f5DHvu39pvYIdOdD42q9zaeb28dP
/QrFLidg2skxLiL3R2ybjbSNES4IIeky4a9rY5LKdCkw85mIRk9T1V80QXOOZI9W1sE9IDuBpMQN
rrRhBeEaCDuHRoyanA6TEclJ7/Wi+z8Z8h0/KC8y6FchMgexOJkEN+UceMdJJGZ0CeuhCFVXOHB0
+2nU9B3oeTu4avfAU+fA7qtHcb+RVIhHnjmNXz+BXkYjlpd9mQ/FFUmmS9GBwhL9PTTVCUwYJWwD
qv6L73n7YDi69Drc/CbC97Gw+YmJtCu3pfztW7VI8hYGKA3xqF0axL+mzXYKp8OBLDWJBFXHGiuo
rW9REUeSoemcZAVdTffOFqNUA2f4hNa/UfBi+ifjk8/XV9yWjIAnVrDU2I5Tsa5q0s9ypo99EWq/
V9GMgcpprU+Blak4yNkQzey//R2hPtSxJRBpW9XXFKFhuvvI4jsAQxoRxMvprhscTrQTnt/iFBk+
Hok/k860l4e9iTeaCa3GVcF+/I7/LbQ6BYR1m/gx8lAFV5WG1ZE/EnVbkOmILfxuQDbjtfLaGviY
XbxArtzj9DFy7k+GOpgnon/5zY3aqmQVMq/DEPIUuSRq5XSqapAiFHb5scl/KY4UVJtftXGoaczQ
OmPZ+x078aI+ePoqeNOi7zE44UiTuJJWGjj+8BgZA3OGQVK+tS0SLz8Ytr1rDW9HTR+0z4zWiPR2
+1Ikw+OnlOj/xw15n6m6PUJvQAhINjamklI1jHvQ9tMeDgQbYlsQtHIBNi0ewVXHJFM05yYHVMe2
O7FoMp/UBFvrQ3CPhbS2Hj3PEgcqMzPUgdRvRTxZ0Y/XSkJJ3GTaCcklYXtBUeZjRiHkY2WA2vjn
d0DxwnfVXU6XQanv7SqYkssfPPs3y5/doJPhKcXpI/FK0+GmX8pd7eS9t/cW+K+RrXVDNn0ttORE
8heMYE9UH+Bd14X6xMTqjIlw3L6cJ0ezf5Qv1bqDaUZj3wSaTZ7niBw6rhi8w9de1RrvZGYPLVUa
5q9l3S9+mzFnD+WxlZwOYa5RelLa7/4LK9HzE4ljTBJBxt6ML5O5+pD6up21NoND+zZblu7bt3fK
/PbY6gCjXzNDKyRhWnchk6pAQB/kGLXd8K+ceV/lCB6c/kiFhBzAVTKezfC3suozTRVv4oQCvBTX
3rkcVFIPKKLSC06SX994LBFcNU575Eh1WsaHCgRDrp4Kh/tuUikabF53vgQpb1IcZi5qDYsI98kE
ByIhuIrvjTMbHtlVvzzN12OlPuDi+xb/QwcYWSxMRS1slYi1uxvx1qal4jDc+1nQIDje0UCp2Q0T
Hg1B4oK3bKCioDYtPIvyrxnEtJ2viFhlJtvV1Jk10p+lL3aWPfOi0DbGiCS9oXCgKJFLmorGKkvF
NzvnHxlurb8Ru0nt9orRwfekLlMOgN5l85Xry3jMRXopGOIXfHqWFhK9OQ8JbnJcKMJ5vpEtOkqi
ooy9n7g0BqOotqn9D7wF0OMrHNRh3hkw9jI9KjYTZn3oa7nP3zLb1J4ksT7v1bCRqZl+a2vubKTI
YrriUtx5NhrELZRAkSR8R/uI/vUtYGICFLomGM/V4N1jBvqPXA9U+EL9sdLiunP7gMPW+Phc7rPI
xyn8tVBPONboteAfK1VolI4LjeHea+ojliOQPr6C64MN9UPf0sJ/HkEi4L4oB+I57UclIFX3fZib
7J14Zn3Dx9Jgc0cvDRud13NxFc5WqRFlYgkTN+Aki9bYEQ4RJNH32ip95mad/W41HVLf9KAKGwaF
1+I6tKN9FRhdsIYTb0Q+T0xhh2os+QPNZaMTwCKvGKY7Ht7Vvb4wEeSjB7Y/hfahk/X40TkhLFF6
0ITzCKykzabmb/z14xu+pKg9qrC2j907+c6p23z0F4RaZMiZhTqBFoGsOyhGwewqw1eZU3YKHBGo
JhsvNu4xIi6yUZYM9oa4cJGr0hxqYW8EaE6/IkueTbNraS8t6mn3tVQxXe6V00t4T0dUPfzqzvxq
OkcMZKFUfB5I/1kGhD8e0RxpI1u9vTv8ZykwoH6nzfOXXnR0ydm6ZiV14C+aVguYqvNJl6d07vpA
smTgT8/uEEjXggq0AM2p6T5rsRax9vsbZRXlTl3i2OI25razmtxHK4Q3Mkhl7fyohTc8CD+7vrp8
pD8kaXaDRLGblmfGDY9Kz1EZJHLn5ekaJ1YUqSTF5zZFu+gqpF3QjMljZrJLgZtshxpNLU0EDKaO
FvhjxN+FenzAVxlKdH/pZU8J+Aep8OMnK9Tlyrj7tvgTZ+gXtG7ATlxFL2R4GpWCr2/ySyoQaC4i
KtymCduWh7vjtwP0AbQTLvchn6utE1lsIh2zK64nYQPXu/hvDDRxeqeuFtIsib0AAu5GmzJjSf5x
YBXmbm497UNQEjfzbuBh794QtxU7MnzOQ2uQxLPnGFEadb/W5oRxRbXGKS6J/GegbFWqCXqOdoor
1WXn5Ub1mRmAE6R38uvQ/HgtwIHZp9UPM/Vm9/BnkFUh98qjhCP8DK4gAU0L7AwR/aDK/8G0KOFy
Wu2X7WScJRZbjcsQumjRDdyM0o3DrIvd6YzaE7Lt73iDKMvTdYn8m1DKFITg0n4HT+e+FnCZBV6b
y2dkps+Jn+fri5G+/q0EbOgwAAFsAZO4GfR21w1i9DW4uFUXRbu9pjXoaj3lcz6QELNf3VokMY36
iBDXuPyRINKgntd3K1LEf63H9ftjoeefU1nQ9f86/m5QdH5S+3gvuwwgpGQoQXkZQ5Yjq+Wtns13
PcZe9WyJlScNZn+xsCB/jPOIEFYpQGKyHcI+GwLbJsNkbLNsAYBmgNX6xbmGuHoUPdAjHYCr9i86
ioIhzifd3+FX/aySUKV3fAYndVfD+puUEbMfJQoGUU+fEni30D5kAugHEtcaVPt+TJX7J4Mg5xl5
dKcFfESVWo5DXwdTDbhGMRzBOZkm7Wp8uVGEQlzAYLN9EWP4zvOF+ZxlaXdiIVHKcxHGxTx2cFir
iBRBryX4xHuw2gNAqLAqV17TUNoSUTEE7W/XJWPmsQjU7VGfnrt54qymE1cL3td5rxBdkxh+UOBI
83u0LL0Oi8rSlvSHri+y6O+5xLe/NzkahIwTLaGDtNlQpcKCErc0CExrJhIH/MtWwcGFlrdjCPdE
bZL5g3E7Gj5cKVVkku3bB+B/7aPHqaaef378Y9hUTjbHu9XyDhaMObktK9BOJ7EnIX5oItuyY1og
QYBWJ/adJfo5PSk5wccp+RaCdjPNrV3Gsg/neud/iljhvAq/iFC4VTTJv119BbO4MD7gJdnguDx6
fchYsi3iwqy1/qHI9QnAiF3jrXda+DZEWxO+o2WHlrS97NHIHW/qhcyi88LzwSpqJeZ4t7lqZNOg
f9zHyw88MxfcifV744UuG1HD7WiE+4PMnxyaTaufQ9szHYgIfJUSdjV3Y+w9lXwyU4jcNjDOIihU
6fRlEmgFWrEmbiJ6uKkA3C2DBsQXrqHxtF/XDLaXMl+UGlHyuF9yX/mec+hKK3ZNluIJfiEishNT
83Wzczk/E22xlV7QsmTfqnZ+512nPCQr8A8NjgORIyAIJih0YLo2kRSgQ3bAPUTjc6oyL5/PumXf
pnUz1AC+FCSWkI36/Ou5aS1Kz+ZeYeAwTtEQTi1SwOIPI/yhAJKQwCZfyRTHKv1HxyrK2HtUA7hb
RaTRxKAAF2UQ9yMrLgA94dX2sszKQJGwoegXMtd92XjoyE6il7OoZ4G5yAo7JgcvvA69mj3NAEIc
nAFS6m6jAFtyEScMiaRHZQI2F2ePYwBmEF58xBVBlp7CsOYH5oWIsta0TpVDF/p8eY0Vh9IIG+13
2m58Hzz1KBPG367iTCkXiFdow2v80fkdux3vDyvGAGVGsABP8XoKRMWotLV+jCAtcLR4LxlgSjb3
KT0W90VaGrRFoURjA1Cy2FJTf5cUMqhStDB90B+4UHhwDSDgVla5G1JUU49ueSeRyz2dJTp8Pne8
TnS0jE7c2YU6xfp8E5em6JiZqOB8y+Gabenf/vlLVBNyYjDOhdUKnc3iz8xzWE2N3NHcsHIbsr7w
cZv5J1/9wLYx8rZpcYNkJy5YcWZ3jc+LJ7GFGbo+MkCoW7MWJzK8fgen5sBHe87YA1P/02l5Fqf7
TjGjNvllmnd/R7ReWke1Hpr/ChZlpJvHb5Bt20GuyKK4zQ8BVUgI3OnZJbAAyd+P8rVBr6htq5oK
n2M4GpcyhhwQ/gabVjc97ldYuZvYMO2Ltkd0RDcRNI4M2BRXDV7tc2q3qlVsm/qnWktVqnN2igvk
XLb5mAMaBVC3e/Q2UdNGVGgY5TyIiQw0WOZ2TuDhnIvO5YFSo/lzu7xroodcdEefJWHKoyyDvwyt
3duP85p8/ACsPmxXeZQrmP4fTv0W590Nru2Gii5UUnu2EpNoIF2HLj32iar2OZYQQX7zcO1O6vCC
H9dStAPcDp/085KOET1b5xrrC9eKqFZmVlIwONGmKdx2vb9wZTZ3IZFDEAhrbMjhdT/mfVYEWC1e
AJWGE9b2iibNswcCGuPLOiZBygnMEPI4IyUOD6bWGaNer7hyGRNoH0WMpEX3WGDtHvuxlkw3wz9D
HXOKPdLlcONS2aeKgi2LA3GF8o4+IaMiVFZfSudcLSUcqCQu3C6d0Y+y3eMNhEkv4GUbC0Vb3lL/
hN+lvbeiNwf5aWusXge4jhv7M8muFt0HKSj5KKHrK3on+GWTFI4dSjlSUdG6gWYT+GvU3+BHIpTJ
yv9Ome7qNIHGpzdGcwXxkDxBzcc4iRvSNQZUTonZ07YwtySAXacGN+fy+keCMNkEcgEHhGPTR446
OEe0ZfPICq1QO4mlVEGpib0VAoKJHFcQELiV6qaItaIhFp4e1gjBEMl7YX7CtPNqA9jfsTZHJeWO
GT0sglvAee22ULZP9n5FfDTHxtK08EIN0Dh/1SIMtDRBZICiUUAeMHHvl5lTjWRUnjIsZgPrrQVE
YzTuRVWVzB+6JSB6K5po6I/IG47Ep6jhIJVmZosG5HnsuanOIn3mDZdnr0LP+4mnAQmIc/+PxNa5
1fWicaxUdlymB+XZ/kTFENbZeEDDhXD59j8AYFOY1cupYZgUEdkrIeOPYhnGkcwpKT5NnX00GJ83
bf+L4336GaHq2quF9Da4NDgzMyRnp+mqPtq7T52ekAzjbM5pUs5dFYFL4no067nMrKmNA6tSlX+1
QBPPChQcEch6fNu7WsQFICcOEx/0mqA5KbIaarui9P3EZdVwdfcHaOKP6XCwXEz3ekzVmE/YLZnV
M+nXbe+Hf8KNOPrmBOjjjI1+4sr6aKtok2F1uosbUQJ+pPnAM/MMug+dImbl/Ay/TjB4GwlqN6RL
TG0UsmmEGnzyMQn2HTFsFpm2qCH1KibBgM4nvPsUu+uNthisXsP87al0skAtIljTExbB06oQyerY
zIk4+FdedyCFQROzHfXJ0q2sJ+q2g2pFn/KO00h0CltWZJ/7yGJYYHg9y+dq+FHouX3Hxo4wQ+se
SAfm5kOBHQwsDh/pRFfV8chhbXKlDYCvVYrPwp7cRLfqq6GLQMJlKdK9b74qR9iTt2lDkmD8Pdnm
wem7FtxYymOhei1aRsXMq+q2TbU05BNRzoO8xCLtKSo7xjfD0KWcwF8OTGa0V/b6j7Q9XHRcJrR9
fRDBE+PMFmJZB92E8k+j7R416qKWrrinzG+0o/9b7wbGZdM7WeSuw4F1zzs3RER4IzeBCc7cZ29e
xi/ZDhsThaNi/dxYoQHdiLREmo4OIbfIfkk8fK2YdUuK7Rznbremy3MAHz0hVQ7UDYGqGZPMO2Wz
3c7AX/LpJH0RCvpBhZIAx/w6Uh7LTSEb5nmdVFupfxYIqzKU0eGWwoIgmaklA6gp+a6cLKkw23jU
t5g7bY6RBLKedQrbOGKzL1DMgxn5vxDnTRsBbNTgh8/KVfC3MLCHwa2LUm6Q+oYTQeylgCV3CdWV
PyRRq2/C5gcxzZ/QirHobwFiDFdE0yM0nhFcZ/GVMWxwG2E77VSQ4XYksv6vnNHw0/CEIimaM0GX
va/N7ys0BZ8Lozos2xKhWEOmO38x8/xCybcc7jMx7SBz9YYXveJeK55ryMCnYNZxZ2rLXYCzWI6C
DSj+hL9Z5XLQELlSdp/K5bKyBLOz5uAMYt9Q7dECkHEsm4w2YAEQ/ISLyyGFKunDhVrbjhlS1dmm
eAemCojhZa2xYfKIXGyK88dYUGWNkzWvDK1RunNW5z0vQXO/ZwNL1vT+2/jTjVribHk2JmC8fZXT
LnbH/GhB4k3xQ3dDBJ6XXKKLj6Z8mCbssy1aqmnviThYk9B5ycqCjfoxBRxGQJEOjxio2GEYQnKQ
JzyWwKKHfTeQ71sDUa2YQ36wnGejNRKxpcZoPiyZb4YTcefeZlxFze7VVvr0FzCpwVQZtWg+Sm1S
hA7vou6BGwLHFeICvcqVtCnFj9MqcBFl1iU0b4AlSRxtbElt9e+NAqxAV5gFIZtFYe9SseY39RXW
KfCHNxPQxLCdKxrWQ+T724o1LUAxazgz+SrqhxlI9lA6vI18VC6Kv2zmH/7LcoxxKwapYFyTwGKy
lNjZ3/wg8JuyoM/8Wkwhfj+Ygj+H+Pqn8wkK0HuOT1Lg09EhXJzTPHF5U995yCa2abY99u9XR1C/
Gaj2GPQBS9VGqbm5zi7fHWy1Cm/Vt7c8AD2xG6oJ1j5T99qnEiXtLt8oF44EUeG0KZgwVViPFfVw
s6tCoNgA9sMK//zvVssTJreDpi7MitoVI+KHCnnaCSv+JF0lJe3DTziTYC2ViqqDpyPswRsN5XRN
nM7jmMVhpDFR0m4rbw3R0sdNiBiSxYxbtjvkRwcjp0VGXVSyjIWqdjYdCHGXPqpQ4uAANx6iaB2W
SSCMvmtpLDkdpqJ1VV2FfLXa+LpYSyc2BDeuieFlF6pDCSWBszJSoIBjJcxJbXkKzEAmf5sZEitl
cjVBJ9Nd9eiAaRpRZaZqv3kKNlBHjZo6tazvH3Da47m7lp+k0hxWcgzv6Cuxd4Z6ATvALPUWAhyy
xPJbWNOggdK0c9kmL6c3vJ/3T4rDc5+m97zSHrrOgMi2V/9JxiTh6xBYAdeeLTHDijBjYjigK083
WK7mzEwQsL03zKryjBXwGN6qOnFP0/8XuG36RNa8cJHY6g4qF+J+keifbYzw8lKqEw19Vuys5A3t
DAOArm7ao2j9S44ugXm4wjWqzCW+U+E1LFuyuGJlidFTmvnnRf7OoDsW/orf2eGH9gvHydj+rd8k
ciOrvdMN8CJDhvhdFx1vb87ymocns/DwtAFGWlBd62i9hKFXAJbs3+/AQU/VhWwESLg77Q465Zyl
7NSjJmsof6Ogp51AwavRBiPk+fio74C7PrKF7IUx2AcgUL1EIZFc6cHlULl3X1qmSmLYUVOVA6M+
Hgn3sqX0511/Y00wRW2qrXY6kLHrCbjs6/rncVB11wzPOlduHZjH3hPYsTauS/uk8gHE955xFS0m
nF1/B5qY4rya8PNmK4ynXcYKvm43DkMc7w0UT9V907xIChorgYP6InnqrFlCCOH5YksHhS2z+rGP
vOB/JzjfFBsoQbaZXI3Su+XzN3J0EDLZEF0tZo6evgX+koi9Rz9Ux0mzESVLjd+p8Sl6HcoQjb1n
KSn+s6IrMbLQmQQv7a7l4Zs8NG4tNwxuwsQdsXWp7u+hdCgFx3kAsYfuVpknnxozbKlA0+d37xBw
RBmOiJeYo2DUf10H70qcx4IERrC3bTsAQrIHHkEOHgGdefWsOALjrhBwzCICEL6gK4T+UzCsqDCz
lofp/9A6RwPogqKLFdwc18aj9yVQdcXIFfkMFysR1egBZqcFgQv32qDdOVrglx9pT1mA0DpPazbx
qrIK3SaAnlPTLtMrZ2uyupM3QcH4Ho5rkh0i//lHXddG0HPFczyBwzhPNZRzFgtmpJc9TVRRwI+Y
wSLK332Awrrt2d3cOcl1rpedaB3bq4gusIwQt72pTfoAoPqH4YqphNYLQ9fSox/+ThG6JN2t9CJy
6IJjNXYSJ/yZX+cAOtepmYEb2i1oooteJiZbcmiOMOFHRsPB9FIPHmz/ex3lZvYAITtqz/Z48lEF
E6CF1bH7CHFfgTaLqp+lTys9hI1HpC+/akA5jOCXKSSkIfkRzTD+7uPdZxBVxNmXA2Ab+ghzXI+S
V8jvTb8426mJvHcqM2aqny+Hg5Nq81ZQj+nShCjT3cM4Y4t3Ac/5weh7v9St8L/JTrIK0JsQC7PJ
2Ce8o67N7fsm3wfAFymDisJYeNRolno5o0WIetpbdgMtUIDeZYvhKaT3z8Ebc+UP9mdpG8Bb+PSy
tzgTTIoTyDLiwLm6JLnNi2AJLVA6lsfGSqeof7NR1OacEdBTuJvqWfoAeV0gPca8WbNX9ga5VhQ0
wJxvz6rrIrnUgSdJFhNNieLSsV80ZdLwlJuq0SYg99WetbCFTDZYKlM5ZzmLl9ZHLz9XD2a0OzTG
I47Jdtk+DVzdfHPNG91ulHIe93SFfj99ZelSiV/09xYUBn1o0aK9vjPIkluHTSb7arbnwJS5Vrvg
BgrVO2GChvJYUBwyyFKG6nLVOKX0EQEbdnYIMT2jFAANm40RJ4DdbDKqxWbeMC3BkvtiRuJACcrV
pdOwwKaVZkC3+YW1xIcCmSB3HQxjk4EQ1TWxE+0WQzjsdr7J5bn5F8NCWMRcGTmTCU/A/OA7DIAJ
h2K02ltqx56H5ClHQyOkksUYrlq7riKKYDOfIEL173kZpyGc5WKmvsNPJsU6fGFrTrmBlv2k4QNk
TMBRvjDseESOejOdqEL83yE51d0AewgiGc1UyVeSe83S7tDiKqFhSkK92+qpHR1yDe+CpajfybAx
Hje3ubpDmFiR1aP/Qgui8WICs6Ytnooogf70h3AmyfqrGliUQVcgWuEZM6F64RbpWun8Xf2325hQ
bB7b6os3y8cmcYtDXAtOcrrJacU4nAPtL4M28WPhaETidAqYHvhUsbEHwWBiepllU3/4Pv1ddpPu
1HIkRkDyJjKryRpmBGs5/nnrWzdRlyQKnI+997cnruSCm8N6h9+66lbeaomRmJZZStmniftwj0OV
6fCSLeQYUf9GJWGABToVJzfDWX3WfWX9KA3DjJ+tlA8XYhkM5WESpRo7qUmoK1wCgQPH2UnqhLgI
bFT/Qb/cVf1/aj1MZ0mqTX6lkbFwgCRJOc4QAzpZLSUKr799KZ7h1TDepGG+awVtxjM7vklsOn9r
IS5TGV/N1hI8c6+3eMdeUwRFJ984SM0pjTYQgiCWVayr+krSyE1UcLzy71OhY3e9yVg60IKPZ4J+
mwBv+4RvjlCmN+pObtMYCE9S+2MYc8XaiI1rOy2wDhfqPCraPaTydSI9hLzta+/ve9FxrVNWzLAe
yKlq7Ouk9AcBLNSXeqhNZ6HIddPgxE+Y5daG22AnMZ34BkSyRraCERlIm0BN0fWfGBknzk+AJtdq
SdxLfui3DBzarQ9ah3wCNY8kSLq6XP4QuhswrPcpCEgVvV78WV4WY+zAu1IniNqnpqlibhwyEsPV
R9ZlikrpMwk0+TPm3Jl4sCZ4cUfAiraUV07TbdsNu9ibJ4olsZ7ybLuU2PBq17SNl4fISFmlgg2B
kbvdTageqgYyKzWfAZIG+JhRO9F4tOuRUYnbx7esMt8cjC6/m18I6nKmbXf5yNOVmARdSGj+gbxh
Fbu5DbEHkQehDbPyVtXZLVvprrCbPWwkOevH5ZLr4oMmV5P13HBoHhdj4hR0PlhFd60bx0VCIAri
VtjSDFe2MkCbXQZ/0n3Ty+lHoIH/1qUON8dGPj7jSLIFG8D2BKgegGWfr3uuefAvMMVsG4n8dTo2
EICUQrV38P9pudhdF/tNMzKYgAlWjYXuyUGjRpi1tGrsQA2BUnCtMCzml1pXyAHYD/vB4que0XVA
B5nHslLF2WEF44ofWTkKV8rPtY8hMJCqxTiUPY6NGRAP1KxVaLT2EwfM854FbnfuPofzEB2fL9PF
xnyhsGxpqkC1z9UsXJKwundGrMXQYVrO91pF+uC6MjqhT2+4cMrwqtBmp+Xz6nVR1pF+xuwsOBgc
SWlB3f+TBtmx+k6V3VLArKNEHHSIlusVAOP4S75N5Y1qnbOmmtYltacmphCA0bgJMaotsoC/GSK9
vvDLMg3E928aEaHFxW/UKUzrYW5qQ+9ZHablRtGW8qao4JHaMvy43PiZ8dZNrFcwms8Y1gISHM02
hsxezepIrytywj/FJmiAfxgKoHddIh51Cc3Le3AUYZiIc+qgpaxUHJvo8vf6/G2qu8XrUYDnukEr
q5po7bUMh6qNRy/AjLvqk3Tr2olEM6epIf1mhqCELhfmzAe9sjyWOQU+f/JiAFFWEakO/uQ/KS5g
F+CXYcK5Uw7mw9jGBabG+nRoLJjZO7sI+mL7XWzTYxaRiqraHQAMa8Jz9/siFA3hL3mdplrgviI7
t9LWnPv0O8nH6A/tHpW6VZCAHZcOPtFP8sRM1sbjGBSghrWcNlzd9UUrQ/lQrxBq00VUbLTyyTLI
N77FTtOOyyFTDbkANNga/F3eUhSDiCPy/oVVcdWMm4ymQgfuidTUPf+rx7f0MWFTkszUVIfsFQrB
NG0yiGBPpyqEKt1tVVyHzWiLLt6LobPlmn3KBGHa9hvY4easAexZyVGXKU5pjlRVSi06naMLw8eg
y8c/+57BGWb4B6HgnZj4vmLhfvY7vRR1AqV3DooqUSlUMRsL/Ivemt8s1rrO0gpyG2A2dVZ/lHf/
aB7wIaWSrCMaD2KtNJQZJXX5uHMmxPCDGuu53Pzor1DD00z9LqiGb+abjkz7Bkw376CX/FF2S0b5
E/2f5MmgkBuBeWFm/zwrYB/AZdJjhapTi39sXXR/MA2GwUVncWeSl+ZVJFA92giTMA2GmI/FZSJk
/QROcIY93nb4tnXrfydIkg20kgd3U8VAiS6Au1CfOYzCYXDoDuberPGjutGsbC6nbgKxoDQ7gkaU
QF5G6qGtaRbvpMfXFFZDPlA66U1eAdYSePK0aMsMtncXv6MLPdhaf77qlEe+XwU1fihP3TGWcVNX
jrFrmfgpHC9ov2DUx0mIZ0ClTxgCfdDMim0yrJ4NzBKhiBmx35nGhvvCIO2qosAL6nxTbzSUlfjb
g1foOQ8xg8vELiTJpXAtPSxvnfNL8wWQ1Wjzbc3ab+oEL/nvvqCUFNsiSmUGlZAa3u2J143yC4K3
DAW0I0RRyGeKy2sjvgFYLxopIarC4ZdGNJfGsxeQi+KAHXN9474SSjeQaY/eabKdIS5tXOoMEXUB
hgvJa6CHZejb+F/g5Q0puT2VLCgSw3NdpAL9J6Te5QRcwcoR1arobfGBaap8kYe6UotlaaSbn9BY
wvukUw6+dXQ15Y+IPC2jIobcf7LZDhJRmSoD101+0IT4u/x2IfLB9aGYAf8Girpy1/4FYgyDc1qr
1db2/j2Y9rXIxe2eopMLFxMFzimIJchff/Hw/BUPet2JGIqgBT1v7UWdzRJEOjFS/4Ntjye45ybm
d8TFdh9IwfzFycl2zDfjIeIG0K2jlSPGRYGyJp/3X31Sy8uhwoTxAdDG06nkj7LwEbu8WABo/qNt
5QRW6f0j6tcDsDMKr007Gs5KAOTz7miBFVYEHTDlWmSPBMDXH9PRoj7xaEruCwKdkC/AOENfan0H
S1uJwFpZsNLeDG/2bPLc5Lpp+9j3EUnfQmxUEnWEM0ClRyrU9z6QzuC0HbU4+wKo3nRHz78ZUuAS
FvrpnDCeflFemU8JgiluiPHW1XTUfatfLL3WTl/cltHInAperJOyF7/orJresiPCHBzFyP25eX6c
d8s40tEunaUAWW1GXHhMwo1ok6L2tX3fRFoVGIcNLKfanKeGY0LGQrnvfnxMzDO3j2PPklm0/Xl6
BCg47IMwJ7gzT9rUGxnNYrLmLZxZGcbZejX11piOuBIOMGssIq2+GW2UIKmWEd/2h4f5IgpGG9oW
HqDFftbG81Z+kf2zMc1amQZV7G7Tw7nOHxpRLpkH42MaLYaCu9beQhRF4TOWmpOwJbsfRW+E9fWt
xVuFySkBv4L2Q8h+N9Jv45+cqMw2jM36fe/4dubdgC0WphmyVkOvs7NEunQbgLJQdCdORRTcMKOC
akVfrvGMWE/wYnMLe71J6RQlLZw+XvAu4LZYfnkZq0/pkhTmudzB7gQUHcXwEx/7XziNOz1WVcwN
Rw/Iad9gyLlVv9PR5VgJ8rG53YGzkCgl2RayzA+kRcLpsRmMrikcF7YLuYovdg5MTmF5ptEqxiNb
zWmHY+H8foD7VLwAx5Is2Udwia3HXEyMzXs8TN/0ceC3PUEi/fn8xLYvpS6ZrRdaF7wV4ZtNXMsY
jjQyWdFRwdbkXoumt7wnEagI7S0eTwfQeyWf35luDIyw5rPmgcpUCpVHez3Hz9GvnE2X2AxzyOwp
4s6svpsHhrxuyk6XL2TfBxZ3uwvQR43WUxzzZuLmZUCWMy2p5qvp/cbDDAGsddiMbMwFCohm8fQz
urbDSbm/VOvggcl4828/5d/0f/wpMMMHJC1Xec85qETunYoaXjhfOzgLpv67tUrsS4BTEqT6Y96L
Az7gpj9hOLUem/gOpX/aOGp2rpOIgN6asM+7wz+v0M62A5XWwQSStAHIjPsQOWraiVJeJh2kNUrn
HlMLsJn8QcZzclHS6kHrhUMNgMY2Qnzn+RzNmgmNTCv9SNq/oMmLwCEbGAkMGWabGrH/MqHAXYpA
Mgn3IsiLWCVRVYjnsfst/n7JTAITVYsmHWyJtjSHj2ZRtDkmfKEKkk5PdHVZz5NIp4HPaFnj+1Ee
uY6vS/Mu6suw69p9nO1sICsMqnkeaoEhfUQPcPsUbNVIWuIX50tutVs2wktTfrqXWG2hoDvlUUNL
+i//7I5cZKEt9jJAVDyyMj60l4V/itCWDj5bSC4f3YIq9M2lU+CaUADXiUruZWJyUdl9wWXQylln
MW/+BdajLilPrzGfcER9kQORfBYO00MtIZmHk9/3QcaVO4mhL8sH2KefpHZYAqK2WJ24Nh6CTru4
esDwERNT/U7m4xb9KTG+OS9Wdx8p33748mUxogiB1nFrGmLch55SVZJU2BJBFN3cNTMxow0zp/ZR
sjU4iGHGCaCg83CYxLrzypQBA2EXVcrRYnPmAuFrBxgXHfJuttVlimn8+yiDwIDuUtFm6eeKpvGO
W712waoZIWdtlxjA1ZSwTX3deFZjsEuBi0eIL6O+XusUCkkBPzBIv7E+TxJx7GTUsJ6tUnT4JBRw
tM2a8505YlKlMHwoGEADEb92o3rb9foGeDazQ1mqMA4NI71D6wpTH2Y7LQIOYFD0bYEE/rbE1MCu
RzvmVBAeT+qSvnmRXMZkDvLjhV2m9wielaLTyht2ZSwRwpQoWWv559QFeIBPWo875tAdiXSB7d4j
ZmsuFLGZcGvofZrhVNhcaGKhAcJhIrZe05sokn/rRLDpQgij7RgQxcOm7te31jbYTWIFXB65pkLF
ZHcbinAkOih/49PaI5d069CHPRhpy+FZfBmKkKrcmJybf0MQLYnaFjTlNYiIxj4bIdGXMLIw0HRN
GnED/DRvF1Lnqnd16GfY9VZwo2zZa0e7ZHhKP1We/WpoxNXxD0kKXXMylKv2hAJ2XM3q78yEzkqm
2SXGKIcGhUUKEjr9wF87t6AFeYoxlv5LvTSrhY7vBd/yWHRL5Mes0lXbdC15YFHR8ESpsFvYQPQw
NAnwQZtQ+kN0Ei6bdMtq0KWZJA5ORu+DUAF4jbqnnxeoEfvaKB8BjhRUJbLEqdZhihL1zQyb5qei
AqieqooGY7BfomjWNcPwSb5fcDQpBBV/0D6Jn4GnFlLnmbzcoQEcoTbDgUsqLddFmmSzg1AFYk1l
4cTQcmnHhhxcUQHXdcGkfuPo8Sy3vUjJUXIWA0W7BUq5blEkResHOTflbtAjIuNOd3q3ca1wCUnz
fOylI2ckz0cKg49g3JqEnP7wYTYbCUX1RJho0a/nT+qWRUx9JSS1vPiNQ7x96HZjbGUY8I22a9fA
HBNPwJhmiRhwWSdYPjUmc0UxhkABf9GcDLIMLFl930VCgttYM9uXnNb3ultmKklsj31ZyJJia36F
q79D+O5/P7dfM9dSt5yEXTmvZTN2kOxVpOzkx/Oumy0dHReE9XJAE8tGv4GabOfR0TG3ys2j6cv/
V+Wad94Q3xAxEa4+Z0dZQzrDzIYNhOIr7SgmsgG7SqyRGLbA3JStNqFOCtmkV9KtoYqbp90DiUvT
31QxFDzKi4HdLDCUG6JMaD5HALvYQYoEgmaQ3Dc/ZmCgw3gpX5KzIyyudTJpJ73yQLQ5+RC/WLih
wI9cWhe/x2gxclwZBT/TG2Jzs+XiqsP4VegGpy8UvNJHwlXofVmPPnSNvNKwfa7V6V8i8OXqqDiw
2HISy2kpJNRcJj0XG1Vhq047zZ4T1XKtJ7pV770d+VoB531yllUKNFELA5mNvoupNDAM6SF0qDNm
UiXY9tLO9W++KCearv5wUC6d/DNtitnwnPado8gcjwHVGb2PsrmRbf0E5lAy8S6bB5LBswZ0QJAy
rkki0W4YbgDeRXbaFRsv/oWFOOehVVEszOfaaphaZQ8ukccD//KoQlnXO69bw/I3RafYnhsQyl0h
asqgZpLSCQcptHvqo2frTQCDvzm2KDbRQUyJ298blXF5tDc/jlvMmW9JwELoL06GH5fvoG6ZUOoz
UJGeJmnVfwXwIXwN1NXHFz8gOW/ij5rfe2sQetH55el/S8ZFjRIAsViKpMAEfiSs270gXissOueQ
nJiWUga8xso7TycRJZwxOOrvaSVgAqWF4KnLI03ozQSruQMETS8OztqW1HSVzZfLHB+15063e1tj
FELXx19AVHQNnQWIc9b/5N4YvLyiU5CrecSGQlgbm9sryro3SHygVJhq01Gw04owvGRAnRs71uoN
VksgAKnz5YLDqySqMZJDSB7bgSmEwVdT3v82s2x8kjr16S3rqsZiM2Y4HjAa2jEz+ewcQ5RXCbsq
ho34NiijfTbOMicCCRjN9JOsoYtpOqAqDolrZsjgnmLGGQPubwlS9dOFP9CkR9uYHCcJRv6xzbHv
Gnqr6ez+PB5ZfvZ5VQoXb2o9CsQtqvpdV48egD0W1C3aXPV+DnmlHt25iLa8obVyY20ZusH+HYUA
0Cur27ko68Dngb84bTe/AXUquQ+ltzHTzDyfNvCLy+gj+zgcwjjRL0YmYuiy3I047k1Eo5iwd2nT
5vwIr9NNlldYFrKmjEr4w0z0CClJMmFF9MOaSbY/EjEHuc6msWaHUXyG1Oh9uSlwD1AZnUetWgky
EtNll6etAFwclIqdodslGD++vTZQd7T5WM4fPBykMERXpN3WU8CiwHoidVh8FonPy3mkoyJyVHrE
ZeVFNF94+t62ATKhizVAbK/2s8AWe5ac+yhM3FR9t70+CIfY5ohkX1IBqlGR/xPNn52QRGUUmXVB
AqIJ6/W1DssRm1IbrGzW6QYsjzB+TBknvoj8Wd6fm7cHLpa6/36apOrEou7mY/60e9CUM44/wChe
/HZXkgGChm65wCnD6sPYgOj8ehBS4WfisbRl9tbRcFAckPKd8SVWUTVJD0aEj8Cegkh0ZLw3l+CK
sUEmpoVDibrOfGzH9P7EudjTHYnIVIzYTP8iDbpp1+MKV315u3KXxIbU08OjwmAsR4GyDgLRf60y
G/EuZDd96MagHt008QvKfch0n7+McjcPvnTe1xShETEDDLxU/TMOEiKdS5d4JBb27L8mCdYLRBh1
eMkSjMbdlOnfcSUsKpB/pW9cruwfET+66887U08FZEs8eEtGgrXTA5y5Q4wOZviOinWlZ1GLa9AV
px/1BgTNLPeyF+n5d0j1SZvAdVr5E6LyTMIDDBAS9HR/ZXrFdvSqeCvdDftwmYmT7mJf8EBoSz7t
DG11t/YH8FAkEZfHGVqv9vqAOAVu4g1OF3w+13n0G+lIXn6JffzMuIDt3RySBMoPPa13fEebWeie
BT6qLf3NGz/37UkTjPnNFJMNbJGZSnRL3511nIa07ZYA8qIF+2gnFFINrW8XoeCB9T6SMXEcrS4s
2dknEZMCwO5wDF98S8O9YIwmw7kaERsKmj2bVa494woPzGyPBhvBQGqFc4gUpGSF6dPSS1kLfQMD
chUDHjU8xt4WEm1eX1XCaa20fR9kql35hq+NP0r7wQDQeEBRtMj8gSNpzvBepLcA8Kabw6Cc7DsX
GkmvYNgOz6oZTjvhn4wUVKazw7ZSxvzJJYO1j4ESmj1aUZqNzslGwjhXx1YzFjPMUssnYl2pyq94
Cl/5wLBrRAp4ATPVM2teLPfRyRJDm1JKm9gEyPuAbKWDIAnkWn3yfTDjSpiCZ8s5ftkPvkD7GYuy
TZCPhHvI5Ot1JGbm4pJ5gzcTA8rdTtrDBe4a3H+DnnhsTro0xzirk1STg/BLOrafQ47LPJ3JkGEa
zqd4r9cK4WuYCOVvhUd7mkXrmk4iaTKH+5OSooR1ajXBE5k5lbYu8JII4ZRkqr/YsR60cQ97InlR
THQO0DK7vBjFrrjeiiWRCl2vz2yleLdH/M8Ta/BkTw7p2t0nG3DGKMTjHKr+tXRgQSZY7/PPnYnN
claqvQHIHaFOYvxVsX+ZC7mSm+Ycs9cIooTa6gmJA60eXaf1ykFyZWmh4V+VEvWVuUJdwvZfQA56
8wm0sDi/p4J6EidLkl+w2tipoRYhHBqwNc57nADgFEWyUqZTvNGc2zsCwoNfcP/D3tamKI+iaHgP
eoMyq3AkBRbaI5fM+y4G02NDG5OiSeO1PKenuJ97AYG3VgLn5dL3lhxVEM+up0Cuf/pR6CGar86G
EJU6tNpBNtZOLt7TBHRpGe3OJDHtMabY2UqwaDH8mKUdOizoG0j/zE8ut9lAJJxzd29G6hymYTmT
3RJURnZJPBR2cenNXsvwpkQLR8AKRxcqGF0qPnZSRU3sRhOMte9+23U+dqEspBKvSuIwc9+Tljyq
KdSNrBSTDVisZv9F4Lus0/7z6VncavoMktHi+oB4DcwUADsw+2sqDe24eCGbfpojtyA0YLCjQo9w
tqkSRgZ9BjY3yUqF8q5J4zpyMLlxsQz3LVVNc0WJDacevPca3gNfYvWIHZ2MKDlYn6G9JGCJ/zH0
XnzT2DPf0M/604JCzJG8u0GkV/jIQcylxrXTD5dGggr5dzKYNviTHFvL3oOA+JgZbWJKLwyrbBAV
JoA1JLTu5dF3oK8qxxJzDJ3Bwme6hmIhfzcsdYOVQTQGTGq4Pe08G8n4RW/o5AbJffJ1dgMOG0yb
+6oSjqrGBIBRL/u1cr6oynGR57/j50COfjfIiBfKSRMvPZpWsgCjc3iJn50Pa1VDRBg8UPjecyi+
9YER43RYFkyHMVWjdKVD182xDp5KT42cJ+rsVePNDmbl90qNtmJkYrfJOAREtMdJCf2QSwotNNIz
UnoAFYmOQQMkIfCuF48EHGtWk6YpSAAAHMBwvNFaxjoYNUqP0+5N2WoQq8kkAmwi+ar4U25tadIg
8bZlUMua1EvTZpXHhchT2WkD6LuzVn05i80KHL1GcrWaU3FOVrflW/LLVnJaGgV1HyklYQGzeGxT
HumfH1lXIbK03D6ggqsLxXtl+ZSWqqvIPf5XETSzmARfq4O8aYxQ3tBFlNKWWv2NwN/ly83y9ieQ
PwEu6rW/V8ykhtMYhyzyAaKrVPedg06OIjwGNtaDDM3mqmUybNwrsDspBWTLAnlNdIjRa3D+UMtB
DELVzhNBBTENJqKS+Yno1bmlg52Yu8A2f66U475XE/BsPqKSc82oj/RYhpuH8US6yoLR+qrit4Td
K5qi8R1RVL3CIke+vWkyq7PTkRq76Daw9e6j7bQrJCvIw+5T4+sDM0Er+cAEEff49ytUCqJcBf0v
Jkm4mNpWJBR48hOf8CYWsZp7L2a87gduqla0JdHqziegd2E7MXmxWveQJXfTAuhkA+HgXRFuEnmV
l5W2Z8aCHvCcHY/vFCblh65aVZcccDiGMpmNVRkDgKf9q2LAZQurKM34ef3USkpFoB5gP+9NA7PH
HyriiKh9I2AcC7CTQ14nbeTbfUQWn0fHcOJkGZo2TzRLNv1WFmsSN2UvDEt5gLimM6CJ6t6DyxKh
GmgUeBQu5oNJip+4cZmTWgwaFJ/bmY90Ss6ZmDBwnFLG1u4d7bTU42kvmVF90Q3jv+oyjusseWBJ
xgwqIFzUjJtqD00ADx074ZdyV80HLCa0ewGHOKsY7KfkLrUTWbdEq1y3l0YexO9Su8glmlmYpPRd
v/UWPsALoqrkFM3IrC8HDZaP99eJPqNrACAE1oVffZ8EfIBXXGhtmbwiX7vNK3P6FceW+E5CCF9n
X/dFEdasEckJ9GBpZmqJaRboeOeFQ8vDM5zScjoVRABl92RNNh+NgHF06i70qK+tMipiHF8+IlAI
mYRFnp/cuBS5g4gIzPn025vOuoJM4x6kuIdDW7JQGQZ/WXzlRV0beWQrThmCLV5YnX3sAVjhog1F
Zvmb8j0L/pHiR/wvPurAFnwq/XfT2e22Ohn/9StuG3R3t5RiozdA+mg0whm/bELi2HWBrSab/aFS
pO5AlmZEDUnayEs8SX1N2YOFCw/f6RykOwjXpbtPEaCcyV8qgr0bXX0+I5+UziwUMMBW16pyuKQ2
SPTVUd54KNjGopqji7Oulgad7OUie5Frf+7aBTFSMF/jGeY8MW9favCZtoYiVAS4h49LjmpzkW7X
Vii2qy4eDks/hXCMu90Wa83hGMJl4JPlG35KmuYFu5QOEWj2y1sJPKi5YpMHk1XpKGPAjKe9q9lE
uAnEP8rvBmC4r+z8E7esrk8mkUOuqb1OIT3dFhYPCR7VZESidc44Ig7qzcDcp48K3JUND/7zZdYz
8CZThbKNc3drW4UsXxZWYMexaI9VwWNtIT9pNjRzhVbbg+U920dvdG33fp8lUFP+JkhsMn2JHAmV
JljbxaRD2lP+ziTqrA8NH2rqyEzc5yTHTBpx21VMubPZYSmXvoPlm9SdpyeeNhEgnol2Vl4NI46Q
+GddIPh3mHlyuh0D2oMS3b9BwjXu9k+T6Z6ZfJZpt2tiN5bhTp8dJEC2QYZNSHX3hG2evPXSZhEg
tJ9mUqTuVFN8WEn+BkCKbFXglA5+fOL6w3FvAEqbXwog+SsHjJdp71/UIqh7a3/LI1ZNtqT2QHGB
/KlvCKslwtLMo61KpWg93HduQ1Ns9EyDYA3s+48mNypxn1oKSZ7fR+CFwNBhUX5S7M0Fi12FoQbX
hntF8MCJZSIjo5u1FSlkpaueQQc0n2XE7/NDk/JfXupuvT4tlaSZyY2dU4SzHERffdiaffohxJIw
/1+OvrvrgLInCnwSfhP9r+kli/ixjGVcwWzAkRz0pl31ReRIgIUNznuFxgS+GvjG6jwS3TtW8TAM
Pn06nP6dTcOBfF3ZS90VjeG/5zCh0j0faINsWnvO9A8/ms/1cF4rfhayWerKBj/trZHciITWbop9
5UUbf09cuBq5UVsqhrjF7Xa+LErDI/skF9A6lahrqG/QfYUTBwBUXLmdr7XKcBb5diWNanZcHFvj
PYhvN8a0hqIjCqRWs8GuIAYo4U3RjcJ2qjGTqPIFVM+5G4JKa/3cvprJWKZB577IYANjLBL+3jMT
VEY3Lpw3DaxkdaVMh4W+ZbcvY1UI18Dvjane4nQfp4vz6jZpamUbcSSXZF7IpA4V2/1r6HHV2lct
+xKyvLs8nVL1CEMmH2N/0dnZ20owPbiMPZBbf0+Np2GvBH8qZZdzLx2HD3efzmWpJjflBBTlsokD
X8fn9YxHj+Y1Apto+XKjhKDgxCKZsAiE3NUyb2krB/lzbcOkw+evWki8bFQhsdsJ1tJwoFmAlx5k
SYJcPv56CZoUcQyac2b6a6eesWD/DoSPvL3o5WCdNlqJef7+HTrm+VFhBkG9LuNVH8RTTSGpIvNe
EZdfNJ6+qT+XN/eG5xR2L7NmlAhbQTVMN6fSVCBx5JhnqcDKcddpbtGMJGol2qFGpVYukmtCAzmN
LYNYFIRzFFDdVNhwQ+EPx1X1uY9o/C2GYtX2NAoVrfnFzWvMYmzm+Kf5aV9bWdyuH2xnnroqJraa
aP1zTQcjPQEwZ/uOLkFv0d6CwMBXG8S9KFcfGKRV+RIE1NeIr55kAbsEfbXiSHFCrJ6e/Y5xE4fC
Mw4s6DiKyCWl92dFAFYhpglYSiOX7nSkkOh6EP2sfPD//sQvOdOawZXa45PLsycs96t8+ACWDPjz
sqq0mdX7YZ4fTDoBuWo0S4cSoasPZVfj/9YGsYuvXG73IAlaI3MD860B38sz/h/4yFzdPfivYa+A
DWC2R+M7bQQYkckBZgrw9AkGe2r7/OeNsoUhvJ3Ry7iJq5Yc+AS/V6behKzab6mXahKFA4+5NDyH
fyeWwcRGqO2YaUv6ytzyUHNQarOjuATb7RQwCxYNSt+nPL9nwg7AvwzYqfTxNxVyeVuxm72py9iB
WNF57FN7J0wqOfvgXxW18nTP5VK3DY5DfG0omDAfVzaaXi1cgqWFG1G1sYBkeoarklSO8OOhjlKa
ZmkV27EOHXB1NpEVdSMA+8Nq7cavhpuid2KYm3cWIwaSmlPOrAn6MocB9Pk4jRWVR+3Mky2x0Hl5
9TxACSFJjFH//BdatJEDLh3ATuTqVNW+sx0NfHatamQerpHYCCPvbnSICSnrj6EY0wwYyVquwfw/
2orH4GYjPaULZ5w+OkjciXdvr5l+po3GVeVU7gDOUninYoRyOk3sTVsflvRD9mn8EhwLOmBTgqsB
ZQ8eJgLhkQ9jmPsTPf/mR7lmGqqpp8ZGtyaAJbah8kGwj1zJGu8Yeil8qMnypfusxcnsbGyXFr/a
FXeXJsxLE6/sojwUak6t3WaqW4nbSNeUQnG0K3SaGd0atdbtXdp6qFX8jgjlOAJ6v9Dfju6meJ8y
3WqG0n1rcqFFdvGRnyf6aQDH92uwlb0Oh6lRN2uteo0zvv4bHGvNUVe38oCz8ntPBKeYJqsCS/aX
hQ+5AwOqV8xVkg0seEQ5cOxczBpiohlfroQguLn+DT202UNpU1laYWZgIcSrm1Xlu3lgmAxBhbqI
HFqot6VUfomFRs25SL3wi2k/U1kgpIFTal6tzq+SqPyecbMz/MilXdAY13fH3W8duzAy6sKREAh3
e/bwyCzjS9CJyM89kA0V63TuKZV4dRhUaiJORnI4kiDWp3XKrH3L7Xi61PXBJAtgbbcNtMg6c9FH
bThPAZ/PqrGCkn3PTzWISpGBpHJUcsxAf5yxXw4JP7OWviA29TyaRtgsXZj24fNWs27DoMxsQZfR
6DEqxxLlFHFnXftkC+If07PkC6MmBzTJJ199KpvgRMgXpgzp5HvYuS/61Z2dP7vuBrvt9uPbUFI0
qjzaKsqazf6hvAHkdPJkdLNE8VRUUl3vf2OzZmX2ADFUee7L0cC+ngBMwJ+IpHvP4oyrkzea+ZrX
j8pmEK5ByON9gDIj+WC0vWulHC3JPau4LfVwSHvBGELBnWwILb1U7+JVowKuJOJl1wLgKHl4zOMw
Lmyom/i2kgTCX94UN7qYjlNKd0DfteDDs2wbAPZcX9bwlY1cFcAkTgUt7s1UMc+SDzubQdfsJpr9
2owO/FDPNAIUtiLPFK7pb9N3oou4c70Ie/EIkwQt6GTizIpdlH0XswLGmul1owvjr5aBBpGAEsIu
k5fqYBKix1YumKVIMhmmNfUI6JTE7h7HovWDPOcya3ggGsJ2bBXg3UJNc+6i+85lWcWEeKCc6bdF
7iMsr8WGsATqDOktH9fFcpiYTsjr+vlzWqprYducz9hRMEjeQ4Ph/qtN/KVmaJfNBUk81o1BwoUt
TzRPlEYwnZko/UbX29AcFTjIAxsjKN8xQPKR2ulIFq8z/XOQwNIa7deIUGZWgW2hlTWSqAvx1kl7
sIUBkl32wg0rZ01Uvqnu7EMS84x+uuxqc4cqb2uozHASyq3iaBW+KSkWLusVa2Hn/8NxGvXk+rtl
S1b6z7gqQdkRvGtPDcGvWjlAYb3qLOadiisUEk0ZU2I5nTC4ttP/+AjNeKFNyUUg75PtsPsR1xlD
4oADgU5QLjg+avqEUj0pqN4vNQ7vgZXBegB7PgvXfTTnS4mZqYzUZYgKa5in48lRGkrOx5C6dSSV
kwrwBP6551NtWmmVQ3sCK97DBRmZag5KC0xNkePx/iPw5FZmI/+cPV2jV9am8KaCekmljmTmInlj
YQ8NFA8RxPzEc/IHnwuczhWl/jlUKubzaU2sp3kIT5YviaCWoO9m0syQA3AUC4oNDHJpseoiykqj
iBOHBEJo7eZD+L50nuElTP4HKN2SCtktzFQZbcM9CsmXg/1TUa5DWVqXosUkpE53gbY89ljeKNt4
sCfYakgEe1jgNttgbQMlEdLadS30V37fqjmZi0+X+CLQResw1zyrxhc8dHOJr7PGwnXPzDkz6VXd
DClDSf9gvcGqyMWledZe8GgjYE9l4q7HalH7EjVHFSN4GXuQNkeHGjH1vGvwoGmF5HvWVfqJ3QiX
gDrGV9ZupY+F9uhTLqgoERsdFHuyPRiAABb9oMQP5IJj6UigYrY+c6AYaPVDKOQcbUmf4QlZCJBd
J7HezaReWx2P/+wwitsqwEmZbcq9YIrjDpyEodiyoT1UP1ilYAo8AwquA1hSQV1AOcTLK+eOET3K
bjwQ+etAhGFAlhgJvAjtQIRGq6z/mkp/z0XrRi9IhlWDqtKviKiu79jHqUHUJ27atNS01B4VFpKU
bcSQj7yBVGbDBmY/EHgwCKoSLGnxyY1NBNiLOQ+h56GGdpQ0JXa/Q6ZWb+nEdvBXVqFrVynJc5pg
ogqyVFU5VRbRQ5EZFJpC/PHGFI1t4xgSmMg/XH+7opxaXCx/zNXCWsyxJzgOx+8LbCuYiB4Pp4/f
cFfQ4jv0jiUInU/FewHlv6kk4rSlO/gFh0i9ZL1V61/ZlkboUHa8yPl7P8xd7Ch3JGq35ql2nNNj
ggQZYdf8O5xyCiFQOT4HbF12vOThN+KZgah0xI5iKAHgMuZTYt6JRrvKH2QSawA5fJ7IqKhTErPV
C16yIU/OiJBsQTG2bSQS707KGg7USodQvvxC+IvNEAtChqzc0LqMLA4n751yRga94Gr1q8PwUQkb
EDe7RsMc8ZgB9Phi+wT3J8J3TsknQ3KVVScujs8EfqW/qwC6whUxtCRGKJqihd85sCu++zXymwcO
Ye0qU452NtTclrR5SlSAY93DAbCPAAld7qxsTylbkc0VgHEe263mJzrEnnRVf/Q4hq/zpX4moV80
gBYyAjcJSgqml/8kh01WHRdCi7wRS+1PcTpZwb+ybsCbmBuYSFhfu0j8bUNgXZkJ8qz62OAhY32t
VcH36O1hxXNc5BLej/aFvfckI2YIkoOlaAyhCMvo9PYwa81r5oUjSgCvmc7kXojnla1hBxa75ypj
ikDvP7EEw4fChof2IHSZnNMNIFNNcnduZbsiYGoOQ/CP1aRorjukNxNXqodCwKlHBPPBQBYYsUk2
JsrH4EwAMC1AY21/9wzGFWOq64LfxjkehO5ejlOtbi/m8uImOrma+e74vYnrawEE/MZ32lwgZ+a/
gBwCNPb/6hU8nAyckITMjrxznQaJef2ZNEW5VV511hzWsnp75VVtirdXfbg0zLXgbBVOujCurhbm
xkcR7aMYa7yZt7TnpBoKz/5pkRZkp59nZ7IMb+mBNHWaLE5v4FPiHXU/PcW1MmaGV5D5IRzFLOBf
MXXesGxc1ZJMnWt6JQwAetZ4Y7j2QhwIfbIGCvSnjJhQeXdPv57s/DxqPueIvQbKzOqlqAiQqZkk
8fwdaZy/I9CYwM+QTROSnccDOjXYn9phYdnehGmayLFGhpMVlKYHsXK+SvP1TFMpn+iBvHbPvo7C
IOSGNtZVRisoSRDcIFf6xE/r2teYFKDXWSRNxhP3Ld6MTR6CL1ypkXfO9pL2cC/eWheIG6DJULcH
9WJNe+BLv4nkm/7tpPDJdk9cmGwI2+Z006ha7GEBmMpo3z78MD+8mBmGQNUY7wVRJ49rT4GQaudd
Bm5n13C5U+nh4bFC0OmFcP9Tr4EokgfUsN7eiXSUjyEfg4/a3Z5y6mugGFsKxcLDgTJfauz/A75e
HRFcIhfa5r8ZQKCe9QOMy0qLmnh0XDIMyZZ13n1p5oj58K6DI6JrSd0o821zoL5eoijvXEf54JJE
Y3WXjjO3fSIgei+p1zcjSGibbGn1CafU0KHCeCE1Y0Ek33Xbs8YcQ+8X7l+yZo3jLJFG6JV/irI9
YoKCe83asECPWCBBWl0TcijUhu2/k7gdymyp5qmvEOEwZJuNU8It9sjXL36m6stZiDsNDpjLQ1fL
NRgyG7vg23iMTdHnlK4LH1vQ/Q3eL9TxaBrPrCsXuYx2X/mUuK5TkVUIeQzB3vQWRymB9QTWrLHZ
M46f6+9CqYEDxBkBDWMxdXRa+Iww1YNjpoXihWP7eH5dCeAdaGuyYLaroy9nPCsXu7ZD+lpMSLb9
VeksuQGW7Iv4bHJTEylEIbli26FtlYwajGvLjy1loyShTmX6oojAFOxYMorUG+a9JV/OIOkT0jpX
y5o3wloObdHkx3PAd7NvaxjzmainAmJX9GZHboLdYQTxms9CBrcCcaF/aDVsZZmDuay9OsKOVT+4
0ULDUlyf9u1yLHmT+sTFG21KfE8imJ4feX5SMczCDsnuqXnTojKAoweWTwc/65MNs4tTk3umxMZE
9zHuRn/KTxlAejgKUkA8Y1qg7T67H46ervs4udqC/i5iijpG37LKHrle0rNkTEMZ3JQ14vojyzKH
e3rEvADuIYUc6gfePaq1QUbyhnHhrOseC9JFCYN5pGMduhm7VRWLpM0iY1mlpclfGkeg1BmipEpV
ZPWu9i7lKMxxzl+dt3/WCqzeiINBkYyOVMtO7seKODzf/3fhsVZla1xf3v5Jik5k0tzeu/6K9biD
l1q9AAofYivudxpjFSmdbyTBld+oq3YTedIp8wC/DuZx1bITNPsupKVFuGkFam+T/8UBrQatSRWM
DHMRLKSEdkFGq9a/BLTvdnPdw6UYSqShFlbGpQPWB92kf8ndAWMYe6tJpZw9fSMd8mE8HiHex0lH
K3lFKSii2xUv4k9ljqvNKvr8MuayoCDOjltfgUvti4IkT3yos6+zodZx8DLntk+8jaV4zBjYIgwe
j/sMsqMt4t2Z0QxfrGebOw9T5kRyWfRJt7hh7ShdCpnlGLWggBRwEh7PvbtyOt/1Bi98dyRW0teF
HscICXtT7lLUfQ6OzJ/BcNcE+4A9ZP4fRT+7LWW+5Toj8guNHCrE5weoqM7z7mbS1TxoNYPelY1w
VPG9huXGpPA011pQCOMB+xO0XcBCdjRAVBjVlogAk7JbgrQFEy1fZ+lj1FBZYruwHpdWvoOq5AQd
wkNu8U6c7kZoRuOrNFeRHZIWT5oTU3mu5AC9CfwR8afQ09PUANa3G0SWGrFpQNVfR/WtQw8XeMlz
N+ueJAwmteV9e6xfqANhg5GwlXtnzf5tM8hi0o/WyYqeHYshO/L5388JBGPZv5tjXNRpONy8n62M
sFEvAnVYwguklcS9LkwyVkyvDfpx2uD8aagskdrj9GMOQEgYwaIfJJupfOR1rJpyAmKTZkY32CCB
r/afP+0RtEvNKEh3jThyIQ3dUymBzNpDuOJ7StXMxB6QpJwbPIVCQ7gAOqxR5TRA8+O1NcJ5kRNC
nxKo5iFoENraKd0GMWk69ScXz/Jua9bP/XGSKzZbX7rq6NJF8RHenw0P3dkx0p1Hfx/ieK5eij3F
JUPOtvRmqDqknajUQvR344rC8HlIVwebscQoeUUTCPc7VcB4Gs4PM80XHrxx3jjOyRQri167Q+WH
0yHjxeuCt2WQFFsadU3RMR2KCACcaUkrBNGljNrDDavytWTrnjiVjfhBv1H1/7ytqFWimsQcV6NB
DDoep70s5bPN4e5bUUBHQEPpoUyDqKEt00nfKOWsoh5f/iS8hyJPEyp/66xjsH9ZXXcalQtBmU5/
rryzGUGbq80SJQfXr590ClzXukt2H4e9TXXlL08+FG6i9eLwl8AvTzoMUkhZR+e/uSPmeHI/9qj2
nHIIUzxRkAwcXEBJ7hikS8jLy6JYE7E4XeMVCrrnKkzD5/xMOCQqyR1aauhv4DWN+IbcKamOBW0U
4WvxxnRMZV+QR8SESA+JEe3fxu6Ig/WRGqwD3Uq5Pbczmq3gr0H4tlC1e5fTOVusAEeND9BNX2H3
CZsKRr/NI4MVMQV0NTEYaS3Nyff/EVXgzbPlXnJK3PGNG8f9PSJuriSJEzucbxVpifKwKkO6BTMI
p8h4c6TvfOA5I+okO0v8wsUMmDWIiwQ4hoIhM+yPdvUeOuICG+oQvPDvzoI6Vx7idv2V/dIMJU1Q
FdOIb02dSJSfdGbAsXTIxDHuIXj4Ihdg29BytXO8/KKR9pAcURdhq2Vo1MEazcZhokNEst9Evisd
I/BP+/sM+kbV0hrpw4OcLu5WsOKN7Z3YfygVsAIj3j6dpY6Cx6wlqlK8QjB0hzxAIJWCF/ZQ1cIL
Vu/1nJVhb9kfO5oXUb/0E/RjbhDH/KgdeIlV1Arlf95bHyzC3JTZoEQ9kNyZmDjnUrOLyUzLtsGN
zGGIeVpkJsE7sUOibTjYWzlF+cyw8bbgaCzxE4ApAxG7GoymFV9/G/+i5h47CvUd6sfOjzaF8IbD
pS77j5zwKkbi9b0tcPHmXPJzHkbRtnIVqj6R8oxKs0VIVe5M1elX+5tiiRm4H91Vdvi4SCTm9pY2
3fvw1UzqQh/Oqkr06SuZPbSsWcf+xAc+zhNTh7s9AoVNgej3MHLv28TlIMN6Lfh0RoRKY8vaOzlc
Q44N3E1l9NhMQTT6Ggxss7SCIpQcBEMMX3uIDBWzlgKXi74Bu5f68OinkL3vurzRaOkVlV9++ymh
GAxJuJnC/UScGin4n94xF82wPfh4NL6vBRW6Vc8gKHpOHK+iDsbCZtJgYyI+N1mTw8wWDGKn+/s1
9aYEfpTtTTB0RaYF/uPn32SO3YBH4cFQLyGAbWqZY3hckeCMASx8R2kavSi+F15js0Et70hFhRe5
t6NKPyJqI4zbWjY5mEh2TlJMPRpBZhHNBvuTAa7zlwnldBJbSGaB79DLDTKALMbIhN1j8SYvBPTf
D1mPhcth4I418Hq+PuO50ijja8CQZ7uWtnFOnz275D/1WyD9svu/eg0eYJ1Mkvox7nyfuG/SClF8
KKdh5akqABw8AUj6sG30PvYZ1GFlzbHX0Vm7gJYXL5F7OOmC3Rc0vTk3163fPWCQ90zdxLtm+fE7
4HWtbzLZb5KkwJWUucy4+KAf8/NZG0cHpjmeVMVDVQuYpRKUGyzYK5U4J2qIHmmrcmlkQ22ig6yx
VTUgGhD++gYo1jQc2F0dFo1WEK3NYQBFEcdkG73zEm4Mws4WpoS1WmJ8H4IJ6XU2Hm1oGxr3dNN4
fPCyvXlh1rH1dElp7/yK1F4qcV7B/f7fC2oGpJ08dNB49sKO7J8ysgmFRYfURdBg4IuzrAd/EQzR
N2JCsVZMFJv2uLccMIV3a4lbHYOifxsy9Boy+WdSBHjvepxq4VWX7UlLteNKKgCjhVP7O4LrF7iA
0Qum3h/WktTspd3HFr68pBTQ20k6lcssg9APVcsnkPDz6/zTIB1liR9acNUBA/VDgTiA0YNmVkWt
3wzlXOCFnA8cmLVBcTQ6HY+nWbDuNCEuEQSJTLr6whZLhhmtQlcEyqQTSMRhG5i+6So0M/7i8ERN
w+WNcnBXO2kTs4Q+XUM8DHF8ruFAQDCcLrn6Qg/4ieRWt1dEcBuvn3C8GRh4CWKhjQpKJ9XFcWAA
lPrbO9XhnAgdb0efBK0vmcDhiZVmyzRAYpniO7hn5mLRsINCty1mCqqJX7GhuOUZZjPxT/g8deKs
nI2Oa1fyY9u8LbgMcQKq4kRRIyxfIpdeq0JKPXrymKDPc1ncsQwcKaLVz/E2idaWnHhs21LCwbbc
JeesZjTTE9nxdatQBQMTlDKipFOVOKwlErh/NmMwn1QdJMqR0wdP/UxdT+Uj8cPB5tUPX7tAOvgO
KJ+8WJ9NmZ9/kCAWXg3v271I/29QIxwXieytIEqa3RkFpkC148G/jE3N1XMrkND75dHjc11XZkGs
LKtryv/wj+Hbrwjrzsndy/kLqOZ4XuygBoFJVceVZqKNwLL6GyktnWN+GR/Ais+hlaNUVq2tqyrx
oNdDfp4UiyPvyfiaCF3Lm7S28QVUJLHu4hNWZudrnFX5M0OjA9T/oNXQEUU64vaxCOuIqgjm/KsF
0Pxi7mpA+PQbnTJgfYwpzYRdsGoihFEaQovNQQc1xyB04uiP3JzUIb1FG1JG7S5U+1BhJe08ujhK
/ID0BrTychiJh8THiwl7OR0CoFHHNI+T3s8mrN9A38xNOOP6LRITgUy2Fq3fvQMT7kZbYcfImBIQ
CAc9SOIHZHzJoK1OHUaRiKE3qUycu7E/O+QcpTw92Ez5ZYpI2H4O6vgFCB8eMsGRB/kQ1FQsWFF1
ppmlKjzofJ7aW5NajsOBBHJiIwbPIBAzOt/2jEIjTzvllQvCaLXOG65C7u4FyZG21ultWkDcLX/l
MIzXpmQY5vcL6z4KWMbzNWO2RV77ht/pupa/jfa5XYc/6anUa4so86/QYm+L1qdf6JpSgGhV+v1t
zf1d1aMyS83I1WoUjFYlirRkgkzwx9qjsvFk8AGGDMSljWwtei5lYGd+ialPJjwUdjdEjU5U4keH
cW5g1wShYuwcJoGmvXXHduOtplyXUxIn38wzKX/0oPEy3BG7LpB6K2RwDQB6r+VnulKpNpC62DuG
v8a67APs0l0Cy8q8NssGMrAi4zNBUKxfQUVMcWUOigpFLKk5JKlWBwdGH7xyEfQ3hLlobmo6ggnW
nYjmJNNfL7e8/pdUQ3LdtpEGqTvD8rHZV7Ijp/CN4KoO7qy6iOc1b/T93dHVccJJokvYYtnQhIOe
t4nvQVN91xu9F1EpEgGg9Evga7iEhMTus/RJFU/L4Q6s+i7q9Uxkc5GjxkuFuZvgafEja4rABaFQ
YgjdLvtfJXs5N0ZSc4wzeIMQLzGY0azfpECivX01j3Jov+CRGZ093NmQUOfWKnbbH60e2ZcnDwbx
r5LWctR+tU4RGJYfirhTrWOXdg1zTsq5G/d9RUOtWJf9/EQmM1FWvHRHdngsM36ZnufpC77jURGU
QJfNbAgQZBRLfsmlLhFx5ehsMpd/IRHXWU6TzxnGeTRKmVmYljfh5gg1uaYzgN5mHhkNjvqE9NJH
iNUIqDxAHb8AljTDSSGbRfV4+0sZ+spOa3yEpWhTZDtt7ImZ2wgw+kqL/IddrvB0nI71oHJdSuyh
qrtxPHpPld4BTIMK1FLKhuT8Be/mkOZ8UbBf4F0YbOp8g7uWCnHvIzU8jA0MPkUGLPIivTzE1g9O
muzRTzWQ+LXov6OjzKIQW1hXzb63TVn60Drxvyy6+IGPwVqp5GbuECMfakwQb2Is4RMa3ZDXybJO
Bp7fH1heVduXOBESkgHGuV/BBRmSggPwn/JGFJSuxVj9EfLUqHYXsLoQ4b5PJmi9ez0K5BZwnOlV
sLgGBJP1RBV9CrRwDtX2T2Tu4Z1cFDfpiWId0XHClv9ffpiDxRlSlxKi5W/lYD4G0Hl3K48bbuIy
8rEZrXsEDXI2YUnMQJc2GZPDCrn7VWkkvMzhnWrCWe4TAn+mWV9dxgvHSo3q8ju/eqPhUwjwJvYP
ZGBgEG1SXV14XP5FjqKtqv37I6+hgpjE5kM9yHFpCnF0SCmfJH2Upbg8y8o5BLMp0iiYyf6/7yQR
aMAR9orVjEBVOHujzWQONulc4SNX65Z0kqDEmm5NYOjkJWu9UFUhSR/o9xBOMjaPa/kjVfgs0UZC
3pn39VT6KwTCG+ShJck6Evh9OYpVcIZgFXwAH2WKN5LLTcOaedJ7yeaIuJXsKWD+hFwisjIc7GsC
vEvdSZF/gpFeNXraarcACjgv/wDyJJ34Wdc2syik8IMloS6A2sHuAu6IJ3OM2HQLJeG/R3CQ0bob
aNJq8iL8GCtKzEyXyxCPO4q1N39E7jQmtFnWOdoaidfqvhI5pqKmhyQfoYyaiGAumCvRT6XL4OQn
STVq2ViAvC+HsLutjNozsOYUSGgMQkMzRirPqWc2RAosqOVvZ2ln/QX03g0lHLGO4E+gxdAhQ3iX
0ZsxHTmBX+epvjz29Mo0CdAffUwtxMbOe7RlBQ0AQceXBeUMa4s1MQYUTlM3uzN6xuHfkBbS5K1M
J7mhrtYfBcc1lEHcZ8x9w0QoqbkUwOOsDy/VmfuZGVmcFo8bb/KTBcW42iRaaM1Tg8VPPbLkM9MN
Ekn0UOjxhqfhqHfa2Zru7T4MUDU9xT6uJIwr4czoGJLpaxtZ8GeFJj8eYcZFzQzkT4rjbZk5lVfz
3duTWgp38A22NU9AMD0HhUq7ljbvYS7epapPiDMpPdeA4j15DC9k8+pyIvXaxLT54yH//otygysV
hkbak3eKhYXbzsD/kHcWWcL2TNnj8BXzB6gnPylKoiOJvQ4r9vcFGX4vq87KwkHyhCk0NPrHXLLV
VVrJoo6y5jOeBmOyYy7jyUGvl15M8yg/wtb7ofgwlTTZw4BJyk6PSD9oLn2TIpmmS5VQWEzMpAOo
hD5gkRNb6R/X7NLvrYcmQnnOKeNG/T6DBtCnTIE5zpnYwAu1da5808QnahUQto3vLB1vTyAbX0Yb
z0JVtfN07dDhpN+uRrMpZxVJZpoNFi/yA1jTHdB9LSpxF5oYMCgTPJN9GtAGRf++MLqcppX41r1j
i1g2pcsONfxnYwzl38Ev6Sk483XuZMeHUgyollIMpSQoPZ2oLvLvIXW/K3vxFKufcY62hSR5NM+k
RgtFoypOWg77qP7iVV7Zx6jAqZYHnpzTokoFsWmnSUoLO2M6Jg1+A8vFkE7a0Ql4PkgJ6maIBq+0
dLppfI3YkFRgYyctmb1qASePO9C/UyPDo8ywnYLBS1riW97C+2RPEmiSU/n8tnqU33E7moCY+iU7
HdbhjybBwMQ4LWzJQgyH9AHqkQTIBfN3MSFgibM9I6RgUbAkqnlFIv1V+QhiiT7vwDXAabn7KHBJ
H2X8O1iOpfXKzA0NLtZsSem/uJF3x+01af5wFIQjsTLJc1Koe0wrut6XkEIkD0J2iBapn7x9KqgS
O6KLVvsGXS+JQth9C6Gq82qWYsDzRe1D4timBfr71qGwrGMCgY3CQ4jJFU5KI6/Ol+r/p7YLxbnP
QjBpbo8eQ40kujmeddWXCVwR4FoRztZ1jvuVLhs8txssLBK5lU4dm60jPqWTaQIvV+vIQH6TkwIU
9fkv8PCT/sHePgrYYamb6dONrlJL0Yn+bKGJim4nMIJOfgn1KsWJFEjUuKaci96918VLe4BGUtZt
uR+ebJFv/LHCvlYVOF0g6WvG/NxTjB4ZG0/T3FcBIn1I+c0aQRqEG5G4r0t3qwTUj2hkzQdU5Orx
tHU0m8B2ST683Uu2RVcS6sjx2idW06zADbFGfpfSYaJ+dQ9b7nN4O9dg3Un58euylgK+ALAUOMKe
SOh8lk7v+CBM/h/jQeWq1gcGeAsRE/5KiL6v7HQYxwv79M6BoiFP85z/K3NEBRXVGjseoiUpBiZd
Frm9d5opg3+2Xr6dxPUvEOAoowCzAlGP3R6b5f+F5AsN5kCH2qJ2XQT2850IIYD6VoRaJaY2kKhJ
U/E2JZGslT4QI2MUjZ0AgBeYoWjkwPTbRUfmwkT+7vmAeCstRNMRE+P4xU9ubAqfyjicWccPi36d
3WrFyd3QsCpkOWH8W2HsNSku1QMJaTenm6jSnoNm3cF56qd/40h4XFmBDP7ubQhbIrs9vktc5Ihe
YTtznCvRNkep961rSpe5w8p0xtKlwzCthMggURdcXqlOzGH2Hr+eppsEW6UhWvhj7jAsqYd+Jiuw
p44kvs3cHkq3XAE7eGi7aNC7C+nO3+G9T4wC2t5/LWkaQ4D0mdFRr7mczDATEMXDEWM2oVuLoy0b
liAbCDAZDcCR+l2hOeenJANXd9zH50r8Bik67auIMVbmZY9bs5iKVWP5cEdUt8Qps/7g1aSpwpGj
PVUw0crS6r0iu6NaD4jL+Hy3RaU7bLopWuM/nEzBZEGmPgyj9Uv5RpiCIs398oCLmtCz+YtsvYSk
7Xzgi3+w8IeHSYOW6m3eylhetlUcJepq5piwKwkNWZi6AmzEq8qPueyT3js6oBeydqvR9nNrVV12
StbACk3ikkLN/ffnepwPlYF4LvQOqJbI5/Ynkf5/NXNaPTv5qweMRZbmAkfTFwtx/+qJf+TF5G6Q
ovGZrlLwC1jhhPEwggN+AdjbAHmW+K8DjqMU/2Px/rwmQYl2nVExA7LhaR0AEsmqpzdYNp8jP+CT
BOL0JIs4vILKj5eDJN3GgoDyZS4E6Nc2cSFeu7rn7TrI4ZhLd/j8UX9DDzBAdXltsr2aOQA/KW9v
nBi2dn8Cely2jg9J39OMgU7I1j0QcDwpeqazPCNOJb7jVltzad23SMtY2IfR6xPBAtOEFAYVzsSj
RY8UMu4WapNAiy7B/GhUiT4buhi1Bqw05WogPRxa3inpbIahiQb73vnLzg7C3+BxNvu6PhllWJoW
EPSPTCUcJ1lDOOKY3A+wNsBU/fLZ6LJg36vEALiK4Ro7rI1H9FrCT3TUCVUPQGUd6m7XtyNOsB/8
94OH69RG5vza0gwxcaQhy4jLMGnMoE1BRU6h6XkFoqOdi3cROjUB7IOP3qZRYY1Hj6Ni5NDaRbYf
EFD64BPb8iUaxSSbjJpP7Eduedks63BpBkcSPT+t6HxgWRv49L46k9ruGFtHbvw41e/f48tKtAAZ
t+0uKxn/U0+5agteK3XKxBG7ytCgMO0n5Pko08ZzqRHUXnGRitkRqJVwREVe8EofAtwnVv+uslvl
+0O2aq8oriaAihje2Q4QcperydSAunhwLct/JWHUPRy433x6Egk5U9FZUIinpQKExjKMRZqd64+S
SsZwa6evznQR/0q/nNeUQaGWHgZ0bTA6hnEKw7i0W6prAwWEHnGfBEI6IE1mwW6H7j/RhQJd1h2z
XyzxhyxElSMX1tyn8EokuNbPpQjtkgWowk6EuALVCzX6sW6n1BxSWIjM2H4XmxlrZpOZRxO8jdGl
aV3IUnnjvcdE1DpTVQG+BQRmfjlhNF1FC4mlFqK5wmWwS5FzRKrBlO7MyvpNltt18EwIL+tFTyk/
yA15NHvx63RAlngJWC6fgdrVEIh91teqbl4RzOfbFNEtlZZ66zxaLixFvROADOGjQJ5jppkSvr3E
ljQspbnKqcSWcP499Rf8Ur4sdZZNQQrkXWsnLgbUJ/6PTIYOczczRZ3zynCSo75DcuaST8FajvXB
+7VHMSJQ+sB3rwcvsL1Semp1BW5W95rcmacJcw+O6cOjeHWluyH4qN3hFfokv8R3Tyuq1wqpNOJd
kXeepFrTClSxnDu9gdX13WhsD4ZR7YGthXTKvyKIsOqTSx7ORw7kW0JuLYGjNtc4H8eodjxQNURo
M9O9TKbfwrlYrtyFRndonSSjEPWuSsSsmYe6R7ouKTkhfUxnV06pzZQ7bJR55TFo+Be32UiwFNQ6
y0QbykPgp29nkrB/lWfGyAJ9rY1KFCi69e5TMf9b/X7+ZQLz7Eh5bK3vkjJNHC8JB3QAAim4C2E7
5rEa9iMhMjcMgLzbaBmBFg+yKblTzoMTb2xV95a4BhBB4IXYLN8BWnA1tDgWJG75nbBwL0o4O06f
DQNx4DXBflAopxGDqCaTDJVAausqIF0PwEAuSB90T7i9spdw3aIlx2ai0hfL/Bt6i37BlHaYQ60C
oZ7bDm6Oh1/LDXIXGh2LwzK/OCvJeDqzenOCr4Ga1aGBbEzYezMzwKNY8tJ1ACT86PSk0znHTxP2
o/PcHEij6ke6H5eyZH8RoH+34FwBrPhF0cOXK88aZTVkc89VSkXEgTCFX1GeRQd/MlVia3M+3ZYz
N4Yt9Ss4Ec4YKxtPzP9TDCdYe+3ljD6gIo7tMChr2/9clAZ6Bh/+TxNFJ7Sh9NHMXZYHFnuqNjnD
PIK3yJEl9IUnMGON3yC+2CTwX/VR1C2ixcny6WelfS/aO09I+EMjqDxlNsTWMH4VCQt3qxRKhyo3
Se3YjlDM1OMSKqm7U3v9UMNTrpqqeVBxLWyzUVW0Ejwj8YgZff/RB7F8txIJ+UHQfuS059Bc3Dsw
7ttp99Y7j8186A9k5qxQQLyunRxaRyu026atau44VvEnzPCmh/ZTBWp3dXiiEJsvPlvJQ10a4Bqu
ZuStI/dBMp6uCXqn5KcOvGpXnEvvuWvEkQ7S2qBJorz8uHC8lC7/fValFF9KY872YBdRt6Jqegk0
vW3TYhlmkdzCU8AM9BUlchkXaBeUiWSVKSYrRpPIneOXyaj3Prrj6uwOx5gEaIk+qzeq/inH95dL
aQU3Gn8EnCC1kttAhgHti0jQuTfnhzk/9/IhPgs24gcXAmoVi81YjmdGIL4jCtElXU+9oBKUrrhs
TmcJgJDqNXnnP34Mm8U16EhN0mjpZp+9/3ygewbQAAfTUOHrt8tAbxzBmq0nCUshmg2nCz7B5xgd
1q/STDeca0cYPVxoGEUg2++iLc7iiGha7GQr5UHNs6OXHPyDvH5GwNPGdiBePn6Vgd6DCWIWkSQZ
ZVpMhkCN254ZU26Oi4Bbw/HswFKtnRG6jqnyq0KO8rP8TTrY1JLNzo9cVDx8GcltfLPMyQ7LJ2Hk
2i6ved/+VWSEFQDEQbeE6yAxQBylwhsCCPf+EOZTshQNyOd/zRNVIPIMjCZMaKRqlnb+OO1gHLd5
qpA9xb0gl+/qd9+OGLi6mS/W0qN5I4elVPa/wLQaZmtS65lYAxqeRf5TcdKiaeirx83ivCBXjIPH
s5a+tiwkCCY43/4JTwEVETEGhFukI+Qbrr9l/RqNN3TXBwBfNwZ1kONhIt6EncCu2AgEF8S3JDKy
lLyimyAB7VAJ8r72XcNJZ8f8Xm0sHdA87pdNz8BqDdr11Bb67Crt/Ax8yN1hGIswNkrtpBFwoy51
EI3GUoWMT7TbZ1xbJVpbVF7RxAYT/mnyd1mf4uUZQrqU74A6Zd/4wPEfOAhLj/KCLLTXskQvy2PS
B/JIdd/825DwWIAcGscR67EC9iixQ7bTPoez6QWZieAzi+EjfViv5WQy/RRIIwN//I4VCYqFkhrm
LMsTNLVEiH7tx446MfIPeICZ+u/gw13GgMFKJjQtldIumEneH/BoKAuues93OBFv731dN44ljz3L
3zV+9TQ3xmRiO9ewX4xFCnl0xYmlKxHvW56bsBBgwH3AmPQN8nPC5ofmr14wy80Z5m5r2sxrHTz1
xIrghvNRJafmkG+2lrT6nejH78KgmJcd+OyLbWgdt6gvVuHjf3Ao/SaZkMz66d+VtysPm4hlTaJ8
HIi/Ky36gV5t1dhdjy5LRW9dBzikUg606L7r29UYf0JloSDK95tHbp9CU6XO9JqXQmJJZOq0U2XK
6YQIfIYbwta15tfSZvjiHIbFNt/no6iOXnpWiI4zryc1jN+Q/B7JNv/nKY9A68fsHhAKYhp8oEdz
Elqp379XLuBmT/vrTmkAct7XqOhdlQ6ROWHay0JVBUAdbTQD0dzOZaQPIKvOqd+/mBlAj6fp/1vD
SXibERjITAuhtSYVx+tQHixlgMmcUOd6vev8AID/bdd+VkT3815UvN2YzQd/dTFFr/ecuNyM2sqM
dcYkYDthgr2JCdG88M4xB1dZBqyCXqGyNptmp/N/ZeRHaOwXvFgId4wKST38Iq6AM/pWp7ccm4nT
7NSJzSwCmC5Zayc7f8etPs/7jre+gPZ66f452d6AK/k+4v3qlqUvdvEhGbTkPCX/pHgNAL6YnRwm
9O9nnhIRTv6lG+HVH6uvm38wIwEh419OmxbyareNO9JLFfiBVeDgzIuALT3/0Kx2ZNmRgOeeAKzN
9uunNcKqFVbiDHvrv+ZktyY8XklV7ObKTQ8Yri+BmvacBpSSQdqkYdhcrkhtM22qKu4VbIIpusk+
GmT4Z7U7tCFpcQRKHjYKRF9KTqAj2nfl+ZBwS0Ieo+yLdwpax74deama1YTK5x5OPVyDtV4XKgIx
p6Pi4e2uD8dZXbZsCKTw+3t1nAaQob/Ub92SPQER8hTJFkZyiyDQ07nKle3MASTXnWI/Vd89dZc+
ARnV8cjhR+nLx8RnD0R9H3cMdel8EPyxG/pT4CTeU3IjIdH4Il7ArJUMp2L0liebQLjJKxPJqf7o
iIWyfT7UK3l4+a5BGswKzT1uc6nUFEygMsaPE/d1SzD/bKkzJlsf3EpjAUMdfEUFdxv4i0PWtBpg
jylTfDs43XgFVl9dux2Ebzn9bK7Q7rjBRLXCUgTIFLnla/piU5lLFnD5fQPv7ba3jzgNcce6iEUb
HF+5OdTFndvMiRnQpQySWxEotQG3YnmSZ/utpE0iUXEWTQAAQ0Xa6HaPh33PZ2Yo4BeCMqCVn3UO
vAmN0uxhpguNPy35rSMCI6HUuvrVJqKTBc97KurgcrPNhgx42uZWrtdcEninfPqKoLyDEVMZ9alC
o9kbdxxgoP/k8C1dNjOJFjhvYXF2hSBPocRzfEiQJ3ASdWsYcHt94cBc3FYHppNWpdwngpwM8mNG
+ZkCbIdzepGb7pz+vPwKH2+vpt2jh+aMewld9MBXmKCSN64mIOzHMlV50W6bIVNyISH2UWhYvoKR
bRZRKX5xoZbZtDrwGfKytobssUcMTnZgriePIRf/5k3fso46UO/PTL+TNtKixk8WpnXz33tPHlHN
5+uGfZ7RSY6QY1efeo7qLslEXumG+r7d1/cpjWxhWimF0k+aPv0XqLsDZA4JomTZnU7p94ancjzX
UqR0KrDm9j8eLXie8fGU6wIBqtslqmbx9cLtkj5iL2ujm/mnbDinqck6VV7HT0fpndoYfYQxqy2h
rS7VWfA8418vEs+hSWTl8o12CGOCGOmKF5NFlykdqg1mRjUn1CjlzOrfF3WxlW54Y77OhyOdy7Ov
xp2dQq4hY85y8z8lKUxokON0/MS2krmlojJiJP7JbQnXks5ipVqFfv+DESRW6aq9kjpjwhvBHoZB
goZDK7Hozed8dT6cEQJkpAE26bkoip95WLArwHK5wPFUIlZaaVGnHo6NgBiO2eNnaRLr66fmu4qy
m6l22AdFmjilmv58eppUmU9RXETuB3yiMhxY2nm0oc3s1lF/q59wpl9G/m2AVWrK2SgQUQ2/Ofme
H7oEkZZx5BAjXvSOKVCW3NiakglHQMIHEGOEXHjQMIeENGV/biYwC6bVmzhP4bfqO9MdC10i9gJC
lhoaps/EJcHVUPNwPXDeLP11p4VvqdaZx0p9TvkRz7sP8o1BwOVkj7V7MxfSnynOfUKKxNmqR+Yr
pnbXr3H71ewztyOpUALifXazizDNT8+g4VuZhwsGvPCe+mZxhHcO0V8mw90pJk2piNVZbL9301T3
tlhphavLKStdunymNPk8BayauF8FWYluCRuKbx2Zw10IHRo2prdhoCdIHtmiGy0CzZSRustdcwBf
Ut2rbr8r8BQ6mPq7yT7lYZZeWh68NSPVJuvgJAy7heEQAT8qZz1vv4ZwhhQUu+rVgUjtn13eHuk/
449Xmu7mcH1Jgxy7dKx1swkGRUKjbcEtEjwEr7yDZv6OdCTaZJ0+zhXs7I5HCG2iMiD40nOg6BtR
GkOacml7aRfc6H8V9cTkHyb02LAIoE/VkanMzqpFA032+X8XNa+5iBcS9MrHbnU/u4l8UxTmjtI2
LF4sKL78Sdo6pgSySzAgsNhvkBXs4Dpz0aRvMdTQv1mD1B8WXRsLiIkpHytYB17MuEWaqOa5pFhd
tLqlJQ8jqC8+m96JDJBCL4KOdDql1bY6iiOb66mcSw4oeUBLW0T4HSZPeCC6HshXFkmKzee87w9E
HUZFvCRpWZaV2qpOkXjYDJ4Be4s1hmIZZUZbpsNFWU8mL4UdFyznAAiPUZ9nRNa1aIv72TNF58MH
skNMdiZeXqFBRHYL7ZCmJ1NrfSifu1LboWrX4oH7APoxVVoQ2t7m7korr/h3C81gCMFpin5O9PdC
1V8FgU3t7CKU6LrCO5XSMTHm4i794mZR9J+ttQZMnQJFuae0Zl/7YX/RL9nfN1IArFFAcjy71b2M
cJsl8JNgJiFa72WoHXANfEF/ZeKsEz6lXFSj5zFR1JmP9R0H1ptN4iuGFxzTOzMNFRg1kW4ofEDm
XI71ey/k1wclUyU9Xa4V8kkOolNDojt4WK5wK6oOLYw5fSN0kcjI1WX020QPyz2md1dmJATzE1oD
AWOdKbl6psFF0O/WRhuib75iEHXN/D5pzks8DwSy1+sMASVTRJ4EPWOq8REj2kESoWhAfWLbl8Xq
Yn+nEGvBFZhpKIyLo32Mr/9VOxdtrd2tkCyM5TIlg7GwO1ODOD34Qriwf/cKp1GWrQBkZuysMdvE
gCPyh9pVadOrU4aEEsE+KNhANw8MUhtnB5WxR6r6sAbZ7FdgAXbtx5AXr9MX4hB8WGqGMJT/4Sh/
MoDiL9Tq5JKuFxp4eUSUGuSKljax6NZNCPElWQQX6DitdvUZZucmZwZzUpk1sf27HZNz3Y/G2Bkf
HIvRBoutgJUO1uwj3Y/YxEItTzU3YnLZJFMdH8fSjn9uOPr1yS+ZB/VZ+LwIxIKOxbZXirUI8r4m
Yx961M5nYa3Fne1/oN2WiJQHBYI6p42cLif1qXlTdiUn6JUSbWftcE8DCxB16uzcPAnWHIEkDwmw
l2F05FT5aruNZKI8aBDzCTPUmF9p2x/cycTpA1SQHKK1FdLfvUoArclj+T2amRpQQyKWCeFduyNe
HRW4JQC7D85EmWJKObUXTsQ59v10+e5a7QcKGDOgli0c7Z6E26Mq2j+M4u8N4jWuH6b7ogVjhY6C
bVBtJCW2h8qXC109j5Sr3idOEH2rkpgLLrYzkGPqWd8kpxgmmDBdLCoV+pwHqARZOe3oDdSKgKPO
7BWpjzejBJgNrCEDYFSxODaYKa7MK+0CfOYv0uK3AM8hir3pvFY2yf+m9aW/O6LQxdNEaiJHQbuN
gMEp8ekSgfrkB/Y+rO3JW3lHvhKj3sTB869YllBiQk23qCz24t6q9wZ3oDIQbKe6srtolUS8XL8X
AApVZTLHOOMghmOqnSJpHKSKmSQm/39ErxMGqjpf0LAcwuCf5AbtoUho7v/4fME90UXDeZAhRwRn
To+0qX8EEm1t/mmvomZvCgfh46P2jGMw70qyqupNTo3vUMDvfvHa9Q20TDyTEmbc9HdcLsurtRcQ
8UGjSFzLgFq97v1C1AU3g8i6vrQxWpkySHrsi1jfGKB+SD3gGk+x6uxiQhKvhXIt+AWkXLsbhHrY
G3apx1MPGXnEw8NSBa8FkwesEPZEL0o0AQsj4wfd8QIZ11MCG9IhKk2rbgbLcobce96aY+fN8ZMP
j13QCrmN95V+lwW+aLi/x496L/quTuoyEUOREpvgq2j617ohUMUwW1nS2X4lmNN+iNGN57MRcG4L
A5MorBRcJZBwxMHTM8L5fwyUytdp0L0mB/QJ/erbPB0mLR3vX/LSSGVPEC46PVeEpt1GgXFkSMCN
CmFXoU6zunc4jcvHaK1MeXVh5MTYuN/CAUJIJaQf92cUI7WO6ySGau38uaYNKuJZzf3q+4OxzTb6
BSaJx3NuBHI7nqN1v54m0NRXG6OwLrmTRdJfituDtk2hjLE6OkjqaBupIO0vtjlJI3vXSDIH5mJn
wSaQBwDliAM1SwJ4/l8NetwoWdx6UtYujBCw5OpI/IKp4QH/+VKspJg80CvUkI0HK3Gogh9OXJZf
eIiaHvfdHjBQO8F+vjC2Q5VfCyh3CkBRgOICOUp7I9cInFfvgGYN9PeNkd9oPxSBiKVVk8nDFV0n
c0gbnqSIWePoPT0FNMN6bLy/LJ+BWDO9cBesZV/zr6aOwiOaFTOnRvQO/8wWehSJi5kjjUNFNvPg
uxmWBbxfOJWZxFgqJPowIf9zYRj7rCedC2CFqV6VBaFUEf1Jt0rRxX9FsSNH2lqbAiMo6KNZKwDa
qDJmRBeQFtmQbG7ke/9FwwonH+YLu9t9PPWkt8EEko1ndP+lfkXmmw2ldouSKZwugNBKgOy2J8Cr
AeTCwk13QJYGeMctWe8BG9+O2yi9pnliq8R7GuPEClkPM5i+nU7ETGj6R3JeYQFwWJPgFGtXfNWg
iyxY5Qf+LunaSYCFl00B1Bw4XAxwypUaC1eyQfENDPFaXzE6BIaxJMkypdI2+qVs+qRQKwEjeeN3
yKuueH/2ROmuex2bpgYM4ZIX41lk1wbA+lV2Ee6+9ka4FZYtYmYIPeRZFMWkSGJV4A5J8JKbu7Bm
pzcAqUDvt2bafTWkgPoZFWDscLKCTmwaRmhR6OBt63A/svaAMhhU0FVeHSZKCoD82oeecrfPw4iG
I4bwpoHt1n/EmntkJk1PXA3UjsUErG26iUufjIYhIMtFkmk5SrELXvzYHVYBScWQunrvZEo4eYHr
kdMyZLxZHteZRVp/wqhmO0EOoqOUR7qKes2biupNN2HmcOvnLXzYjSGp9P3HgSctFFYzwDLNJ3zL
zh/530h6nkBUdIsB/l05k19GF9LTDowE6kXGTY+/2EIIPRXfAwGtmY8gIecjptqHOb2wBFSDb0uZ
1R51i++PSXWEUTQrytXa2sk4qW2AXjoM/TMgkRMXfS0cHj8a/SLC3KeRO72+lyCuoZ6YsarEjF03
BC2GB4kX25QR+MjgH8mQmQdbR7qxQ/M6heY64DL9yUxrdMO2ri2VOIQojzkMVJIEli2ZYcxhw92L
/fOEg9gAqpohZVYMWzYth0pninW8twt/ZuYz+m/eIwrgNrEaqJGKr1CvZLgpyiC3BYLPmTNmzJDZ
OnpBz3VpaOIrD85IU0G5A6i2nsZU9Ht34oWShAQc0KCRE0K2DYdomgTDWSUODcWEI89kK0k6fFPf
sX78AvSIphpKeZ+ys2rViETl3vQLwQ3WkBB6tyIvZIKeta7anLR3MK61zEa04T1n105FhDzkNvmY
gi1C/hFNlRwq6/3yLMubGOzz/EFoMKe56o4KhmktO1eTqw8hHN8AJP2VTvzrTcMax19abPEOpiC9
9cLJURtkVbVopvrugiomXyY8H7IlQiumJV1nwkXMAj1rOF6404kkZCQDxrhCRy/fm8q0740jnK7r
1ejZw6LS8mGkXUuMOk1z6DG+MSnqc9jYKgapcRdf71YD/dXynxD5dPKBNneurICnhaA8FROBOpqW
jbZZ7mTZGglCJC74+G2pL7vK2xMAb7cR/UV+xytVmGP0OKr4kzL9EL/hGsz2vD9lIWdu2BcBcl+8
gyq+kk/4CcJWaSANJcvACSil8NOpWgUuPkEHledtnurlWlB5oH7/zYemulgLJHvlx5s/g40OPhcr
shr5rlgOKZdrItjy5Mc798FeqtpDeb93ZbEXMlxSfHvktqpFZdrAvRkCU9cYLEoPGcbMS34SXfic
9k1p1zyLJ5j8536VH+5OXewSJ83L0JvVogN0n+vppt8mkp1ZkG2Y5TxbU5RGJUc/uSrLymRoGz9j
87xqYhkEhU85C0LFP4D5O7oJEgv2d51ZPrLxYNS9ILpY8ZVADgT9BOmxrFbvbcucfgZbjXhjeAS9
wUmOgYe4WLmbNYXP8HddFaeiddQWglc39fxfDj/lOC/c+bPes/bR597q/paXcXyl/fgsQ7DiK4mk
PLrvrRf+Q6VxjMYJt/EYdIuJsSbxHSmW4CvjDNdPliRwjUeQh3cDghfXdZn+C2SdTQl9Cc0WVApo
iQpeDdiGbp1pLLkzY+yfdjqH1oMssDDWPTEE6wJz6ZN3BkxrNK2gsqVpzznqJ3bqDg3WybeLmkGi
4ZOnnYAjfTHUdfneqbP43+d8JsLWhWRu4OJGBFM1drNteWgZtPVJchq9Ej9sZ//XAIqOmf4JJQns
EjbyuVXkXlbhWLe9Mu6pQDWuq9TgrWKA4cWRkxjjmRhX0jVuKSG6Gv6J+WXOKwzyLzJo/YzJ+ic2
IkMVI+QGUKj+/4XzkPQoRCPhac2rc0AIeh2KphzarCSD2U6Y01FI97hQOUr/A6Dz0YiL3M6rNyeF
xVyjNZC7D52Rh9K3OYYW4DlzYC1/JyBH78UKbdU1E6XvlAY3pbFiedVSQZYcx3FZzAhRKzOwd4kt
IHrGKsQ7XcD9ry7odhZEJmHVZyAQ50Z9BpcbepaCvj9T8PB8fGwXx6gR4Jc9hthzQFukpcBxVyqx
WHSGLMM1VBfPofXbfLVNltsbQ7DrsSjHpiwqSpHNzSJHcIhpqOWm3vJQmQHrln8tXI52ZVxAcptw
yHxMm65rqWknCBDQCVqLNlYt/5TK23BJ+6R25bzyWxPmNAvMt3ote6ys/rP5ei6WcFj+1qQFdFRV
R1lGfEGeZBGJmy+9DCaa4h8Qt3YfFMA/9wJpNnheSkF9BQUZRrpGqmYNbUBz+YRuxsaF17igbIFi
EozbWVOtObc62qIwsejdkBX73HtginMWEgIJ0HZPpwS2E+Q0CtNmYn2nAMGfxuMxM3GJiNYnJryL
2k17zYe8EXBEJUOcloSASEMUx1MvWXNVfi8g3qtbXcMhhUz4IfhZRahaXKRxgj09uJA+l1Ij+M96
Z+VKkHav5weUbokXBtSZ1c2e2Lgh5XLFRCue/pjiZLp5uuwF5Wy6p4L3qIB3wUeknIMFZfvxhukF
clZ4GO99bQffhfocTi9H22hrRqHtVr2W1dsnWIlAM7FdF8D1Yf1jf/g6bY+jTwOp+ybTaTjxxhPK
dn8DYiNDIej0tt3WHqKxqlC+F9RlCN6fmaV5XSYj7ZVFTuVGueX8ioEls2Zl7cUfbP2odQdUgxVU
AWieO5BLlJF7HDHX8neMecUneZyPfWP54z5gJX01crDfDTBGe5akp0rN+p8qOcyPhRpBQy9MKZCO
nyWZLMvpH5NuMUGeqsGWbFeQKXk02+bgesiHdpG5IpDBZF9GWNhuFckZxyR1z5op1RAvZszOidRv
Rn7foplWtKsavO49QtGQY5FIRSwgPwrA2IUOrAVvZ6F8aXib/8WIriPPIGsxcX8Yqupv2uNeUj48
tlD1bxaIwowB3rzc+onkTN4Vz8USAZgkKjYbaV6SCCEHrMq1K21VdY+AQgfcbc4OIVwdxYDJg9Ga
CWzSen3YesgAv4nMux4Bbm5i+0OPgLFNLbG3oYxY7HoNVMrsKQG1Oaq/ywwrteuhYJhWM3Ajjxf8
j+QE/eYgoEAhnl9Rhog2nsHNnZymDO22Uw9j8vOyAFub7huDwb7OIPURLEK5fuxgUEWKs6EyyCCV
5Ax+94qNHZCp/cl5zhuW5/MAXt9tkMQYAISH3cNXSF72PzhATJ7YVg2XFX9eDo3exFTeEVSVVF3G
wyrHAeGqpAY/olpUUOty0QIYduOLJAFsgndV/+h+aFegZUf1r2gBvNFGuKYhkUKtBr08bfXhVfAa
vICq4DZsxWyLlWPJhYYVws9/f8Jc2Gw9RpQedadT/oeeDtv7GQXFRLcmGpEsbo5Kr/U4SIxwcq16
C+GvRkUfoerzC0VqO9e7uLFVfpXCyU305LpEu/tCBY1SMO6FVMUi806yguJfV/spOQuujtJNlfNZ
vQj0ozVorIWOmcg8ZksSd+psdDow8lUQMNgkQQT/IcIyeb4dFyygpURI9AlUYoyjl8tE7tSVMkRU
F5lLXSvzMbtzE5VZrjvxg8evZtu/xpsvKp3fIIvRO0Az6t92fvKQ0IRLrgqqpLTqTLZil2lUXlI+
OIf+0lZTT09YubBPm4zJuLTXihdxvR9+ZC3JCpQ0Ia1tAlhvqt+pyDJEJkES5ek/cMf1aTbdgRxD
PUNH8pBQo75KZvepGPDdL4ELmAH6FuZmCVJ+zTmn/zwnnLl75muhz0otE9ucdPhf/yLP5xTtBjVx
87Co7h/RC1wY1uIvC6CjjMAYTquiLIOGi3txAMgEJOzWFbq+lCVVEJhWZZlJ3Si2hPOXfTMBn8pO
XuP3Hhtovw==
`pragma protect end_protected
